library verilog;
use verilog.vl_types.all;
entity alu_hier_bench is
end alu_hier_bench;
