
module pfa_95 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n2;

  INVX1 U1 ( .A(Cin), .Y(n2) );
  XOR2X1 U2 ( .A(A), .B(B), .Y(P) );
  AND2X2 U3 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U4 ( .A(P), .B(n2), .Y(S) );
endmodule


module pfa_94 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n2;

  INVX1 U1 ( .A(B), .Y(n1) );
  AND2X2 U2 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U3 ( .A(A), .B(n1), .Y(P) );
  XNOR2X1 U4 ( .A(A), .B(n1), .Y(n2) );
  XOR2X1 U5 ( .A(Cin), .B(n2), .Y(S) );
endmodule


module pfa_93 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n2, n3, n4;

  INVX1 U1 ( .A(B), .Y(n3) );
  INVX1 U2 ( .A(A), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(n2) );
  AND2X2 U4 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U5 ( .A(A), .B(n3), .Y(P) );
  XNOR2X1 U6 ( .A(n2), .B(n3), .Y(n4) );
  XOR2X1 U7 ( .A(Cin), .B(n4), .Y(S) );
endmodule


module pfa_92 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U2 ( .A(A), .B(B), .Y(n1) );
  INVX2 U3 ( .A(n1), .Y(P) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_91 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U2 ( .A(A), .B(B), .Y(n1) );
  INVX2 U3 ( .A(n1), .Y(P) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_90 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  XNOR2X1 U1 ( .A(A), .B(B), .Y(n1) );
  INVX4 U2 ( .A(n1), .Y(P) );
  AND2X2 U3 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_89 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  XNOR2X1 U1 ( .A(Cin), .B(n1), .Y(S) );
  INVX1 U2 ( .A(n1), .Y(P) );
  AND2X2 U3 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U4 ( .A(A), .B(B), .Y(n1) );
endmodule


module pfa_88 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  INVX1 U1 ( .A(n1), .Y(P) );
  AND2X2 U2 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U3 ( .A(A), .B(B), .Y(n1) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_87 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U2 ( .A(A), .B(B), .Y(n1) );
  INVX2 U3 ( .A(n1), .Y(P) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_86 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  INVX1 U2 ( .A(n1), .Y(P) );
  XNOR2X1 U3 ( .A(A), .B(B), .Y(n1) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_85 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n4;

  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  INVX2 U2 ( .A(n4), .Y(P) );
  INVX1 U3 ( .A(n1), .Y(S) );
  XNOR2X1 U4 ( .A(Cin), .B(P), .Y(n1) );
  XNOR2X1 U5 ( .A(A), .B(B), .Y(n4) );
endmodule


module pfa_84 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(A), .B(B), .Y(P) );
  XOR2X1 U3 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_83 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module pfa_82 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module pfa_81 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(A), .B(B), .Y(P) );
  XOR2X1 U3 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_80 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module pfa_79 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n2;

  INVX1 U1 ( .A(Cin), .Y(n2) );
  AND2X2 U2 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U3 ( .A(A), .B(B), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(P) );
  XNOR2X1 U5 ( .A(P), .B(n2), .Y(S) );
endmodule


module pfa_78 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n2, n3;

  INVX1 U1 ( .A(B), .Y(n3) );
  BUFX2 U2 ( .A(n2), .Y(n1) );
  BUFX2 U3 ( .A(A), .Y(n2) );
  AND2X2 U4 ( .A(n2), .B(B), .Y(G) );
  XNOR2X1 U5 ( .A(A), .B(n3), .Y(P) );
  FAX1 U6 ( .A(n1), .B(Cin), .C(B), .YC(), .YS(S) );
endmodule


module pfa_77 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U2 ( .A(A), .B(B), .Y(n1) );
  INVX2 U3 ( .A(n1), .Y(P) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_76 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U2 ( .A(A), .B(B), .Y(n1) );
  INVX2 U3 ( .A(n1), .Y(P) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_75 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U1 ( .A(A), .B(B), .Y(P) );
  AND2X2 U2 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U3 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_74 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U1 ( .A(A), .B(B), .Y(P) );
  AND2X2 U2 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U3 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_73 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U2 ( .A(A), .B(B), .Y(n1) );
  INVX2 U3 ( .A(n1), .Y(P) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_72 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U2 ( .A(Cin), .B(n1), .Y(S) );
  INVX1 U3 ( .A(n1), .Y(P) );
  XNOR2X1 U4 ( .A(A), .B(B), .Y(n1) );
endmodule


module pfa_71 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U2 ( .A(A), .B(B), .Y(n1) );
  INVX2 U3 ( .A(n1), .Y(P) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_70 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(A), .B(B), .Y(P) );
  XOR2X1 U3 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_69 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(A), .B(B), .Y(P) );
  XOR2X1 U3 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_68 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(A), .B(B), .Y(P) );
  XOR2X1 U3 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_67 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module pfa_66 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module pfa_65 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module pfa_64 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module pfa_63 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
endmodule


module pfa_62 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
endmodule


module pfa_61 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U2 ( .A(A), .B(B), .Y(n1) );
  INVX2 U3 ( .A(n1), .Y(P) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_60 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(A), .B(B), .Y(P) );
  XOR2X1 U3 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_59 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U2 ( .A(A), .B(B), .Y(n1) );
  INVX2 U3 ( .A(n1), .Y(P) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_58 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n2, n3;

  XOR2X1 U1 ( .A(A), .B(B), .Y(P) );
  INVX1 U2 ( .A(A), .Y(n2) );
  INVX1 U3 ( .A(n2), .Y(n3) );
  AND2X2 U4 ( .A(n3), .B(B), .Y(G) );
  XOR2X1 U5 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_57 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n2;

  INVX1 U1 ( .A(B), .Y(n2) );
  XNOR2X1 U2 ( .A(A), .B(n2), .Y(P) );
  AND2X2 U3 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_56 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n3, n4;

  AND2X1 U1 ( .A(n4), .B(B), .Y(G) );
  INVX1 U2 ( .A(B), .Y(n3) );
  BUFX2 U3 ( .A(P), .Y(n1) );
  XNOR2X1 U4 ( .A(A), .B(n3), .Y(P) );
  BUFX2 U5 ( .A(A), .Y(n4) );
  XOR2X1 U6 ( .A(Cin), .B(n1), .Y(S) );
endmodule


module pfa_55 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U2 ( .A(A), .B(B), .Y(n1) );
  INVX2 U3 ( .A(n1), .Y(P) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_54 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n3;

  INVX1 U1 ( .A(B), .Y(n3) );
  BUFX2 U2 ( .A(P), .Y(n1) );
  XNOR2X1 U3 ( .A(A), .B(n3), .Y(P) );
  AND2X2 U4 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U5 ( .A(Cin), .B(n1), .Y(S) );
endmodule


module pfa_53 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U1 ( .A(A), .B(B), .Y(P) );
  AND2X2 U2 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U3 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_52 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n2, n4;

  AND2X1 U1 ( .A(n1), .B(B), .Y(G) );
  INVX1 U2 ( .A(B), .Y(n4) );
  BUFX2 U3 ( .A(A), .Y(n1) );
  BUFX2 U4 ( .A(P), .Y(n2) );
  XNOR2X1 U5 ( .A(A), .B(n4), .Y(P) );
  XOR2X1 U6 ( .A(Cin), .B(n2), .Y(S) );
endmodule


module pfa_51 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U2 ( .A(A), .B(B), .Y(n1) );
  INVX2 U3 ( .A(n1), .Y(P) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_50 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  INVX1 U2 ( .A(n1), .Y(P) );
  XNOR2X1 U3 ( .A(A), .B(B), .Y(n1) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_49 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n2;

  AND2X1 U1 ( .A(n1), .B(B), .Y(G) );
  INVX1 U2 ( .A(n2), .Y(P) );
  BUFX2 U3 ( .A(A), .Y(n1) );
  XNOR2X1 U4 ( .A(A), .B(B), .Y(n2) );
  XOR2X1 U5 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_48 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(A), .B(B), .Y(P) );
  XOR2X1 U3 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_47 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
endmodule


module pfa_46 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U2 ( .A(A), .B(B), .Y(n1) );
  INVX2 U3 ( .A(n1), .Y(P) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_45 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U2 ( .A(A), .B(B), .Y(n1) );
  INVX2 U3 ( .A(n1), .Y(P) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_44 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(A), .B(B), .Y(P) );
  XOR2X1 U3 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_43 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U2 ( .A(A), .B(B), .Y(n1) );
  INVX2 U3 ( .A(n1), .Y(P) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_42 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U1 ( .A(A), .B(B), .Y(P) );
  AND2X2 U2 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U3 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_41 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n3;

  INVX1 U1 ( .A(B), .Y(n3) );
  BUFX2 U2 ( .A(P), .Y(n1) );
  XNOR2X1 U3 ( .A(A), .B(n3), .Y(P) );
  AND2X2 U4 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U5 ( .A(Cin), .B(n1), .Y(S) );
endmodule


module pfa_40 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n3;

  INVX1 U1 ( .A(B), .Y(n3) );
  BUFX2 U2 ( .A(P), .Y(n1) );
  XNOR2X1 U3 ( .A(A), .B(n3), .Y(P) );
  AND2X2 U4 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U5 ( .A(Cin), .B(n1), .Y(S) );
endmodule


module pfa_39 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U2 ( .A(A), .B(B), .Y(n1) );
  INVX2 U3 ( .A(n1), .Y(P) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_38 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n3;

  INVX1 U1 ( .A(B), .Y(n3) );
  BUFX2 U2 ( .A(P), .Y(n1) );
  XNOR2X1 U3 ( .A(A), .B(n3), .Y(P) );
  AND2X2 U4 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U5 ( .A(Cin), .B(n1), .Y(S) );
endmodule


module pfa_37 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n2;

  INVX1 U1 ( .A(B), .Y(n2) );
  XNOR2X1 U2 ( .A(A), .B(n2), .Y(P) );
  AND2X2 U3 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_36 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n2, n4;

  XNOR2X1 U1 ( .A(Cin), .B(n1), .Y(S) );
  INVX8 U2 ( .A(n2), .Y(n1) );
  INVX1 U3 ( .A(B), .Y(n4) );
  BUFX2 U4 ( .A(P), .Y(n2) );
  XNOR2X1 U5 ( .A(A), .B(n4), .Y(P) );
  AND2X2 U6 ( .A(A), .B(B), .Y(G) );
endmodule


module pfa_35 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U2 ( .A(Cin), .B(n1), .Y(S) );
  INVX1 U3 ( .A(n1), .Y(P) );
  XNOR2X1 U4 ( .A(A), .B(B), .Y(n1) );
endmodule


module pfa_34 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(A), .B(B), .Y(P) );
  XOR2X1 U3 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_33 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U2 ( .A(Cin), .B(n1), .Y(S) );
  INVX2 U3 ( .A(n1), .Y(P) );
  XNOR2X1 U4 ( .A(A), .B(B), .Y(n1) );
endmodule


module pfa_32 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U2 ( .A(Cin), .B(n1), .Y(S) );
  INVX1 U3 ( .A(n1), .Y(P) );
  XNOR2X1 U4 ( .A(A), .B(B), .Y(n1) );
endmodule


module pfa_31 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n2;

  INVX1 U1 ( .A(Cin), .Y(n2) );
  INVX1 U2 ( .A(n1), .Y(P) );
  AND2X2 U3 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U4 ( .A(A), .B(B), .Y(n1) );
  XNOR2X1 U5 ( .A(P), .B(n2), .Y(S) );
endmodule


module pfa_30 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n3, n4, n5, n6, n7, n8, n9;

  AND2X2 U1 ( .A(A), .B(n9), .Y(n5) );
  AND2X1 U2 ( .A(n7), .B(n8), .Y(n3) );
  INVX1 U3 ( .A(B), .Y(n9) );
  AND2X2 U4 ( .A(n6), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(P) );
  INVX1 U6 ( .A(n3), .Y(n4) );
  INVX1 U7 ( .A(n5), .Y(n6) );
  INVX1 U8 ( .A(A), .Y(n7) );
  INVX1 U9 ( .A(n9), .Y(n8) );
  AND2X2 U10 ( .A(A), .B(B), .Y(G) );
  FAX1 U11 ( .A(A), .B(Cin), .C(B), .YC(), .YS(S) );
endmodule


module pfa_29 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n3, n2;

  INVX1 U1 ( .A(n2), .Y(P) );
  INVX1 U2 ( .A(n2), .Y(n3) );
  AND2X2 U3 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U4 ( .A(A), .B(B), .Y(n2) );
  XOR2X1 U5 ( .A(Cin), .B(n3), .Y(S) );
endmodule


module pfa_28 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n2;

  XOR2X1 U1 ( .A(A), .B(B), .Y(P) );
  BUFX2 U2 ( .A(A), .Y(n2) );
  AND2X2 U3 ( .A(n2), .B(B), .Y(G) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_27 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U2 ( .A(A), .B(B), .Y(n1) );
  INVX2 U3 ( .A(n1), .Y(P) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_26 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U2 ( .A(A), .B(B), .Y(n1) );
  INVX2 U3 ( .A(n1), .Y(P) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_25 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n2;

  AND2X1 U1 ( .A(n1), .B(B), .Y(G) );
  BUFX2 U2 ( .A(A), .Y(n1) );
  XNOR2X1 U3 ( .A(Cin), .B(n2), .Y(S) );
  INVX1 U4 ( .A(n2), .Y(P) );
  XNOR2X1 U5 ( .A(A), .B(B), .Y(n2) );
endmodule


module pfa_24 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n2;

  INVX1 U1 ( .A(P), .Y(n1) );
  XNOR2X1 U2 ( .A(Cin), .B(n1), .Y(S) );
  AND2X2 U3 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U4 ( .A(A), .B(B), .Y(n2) );
  INVX2 U5 ( .A(n2), .Y(P) );
endmodule


module pfa_23 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U2 ( .A(A), .B(B), .Y(n1) );
  INVX2 U3 ( .A(n1), .Y(P) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module pfa_22 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n2, n3, n4, n5;

  XNOR2X1 U1 ( .A(n3), .B(B), .Y(P) );
  INVX1 U2 ( .A(P), .Y(n5) );
  BUFX2 U3 ( .A(Cin), .Y(n2) );
  INVX1 U4 ( .A(A), .Y(n3) );
  INVX1 U5 ( .A(n3), .Y(n4) );
  XNOR2X1 U6 ( .A(n2), .B(n5), .Y(S) );
  AND2X2 U7 ( .A(n4), .B(B), .Y(G) );
endmodule


module pfa_21 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  XNOR2X1 U1 ( .A(Cin), .B(n1), .Y(S) );
  INVX1 U2 ( .A(n1), .Y(P) );
  AND2X2 U3 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U4 ( .A(A), .B(B), .Y(n1) );
endmodule


module pfa_20 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  XOR2X1 U1 ( .A(Cin), .B(P), .Y(S) );
  INVX1 U2 ( .A(n1), .Y(P) );
  AND2X2 U3 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U4 ( .A(A), .B(B), .Y(n1) );
endmodule


module pfa_19 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U2 ( .A(Cin), .B(n1), .Y(S) );
  INVX1 U3 ( .A(n1), .Y(P) );
  XNOR2X1 U4 ( .A(A), .B(B), .Y(n1) );
endmodule


module pfa_18 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U2 ( .A(Cin), .B(n1), .Y(S) );
  INVX1 U3 ( .A(n1), .Y(P) );
  XNOR2X1 U4 ( .A(A), .B(B), .Y(n1) );
endmodule


module pfa_17 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U2 ( .A(Cin), .B(n1), .Y(S) );
  INVX1 U3 ( .A(n1), .Y(P) );
  XNOR2X1 U4 ( .A(A), .B(B), .Y(n1) );
endmodule


module pfa_16 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U2 ( .A(Cin), .B(n1), .Y(S) );
  INVX1 U3 ( .A(n1), .Y(P) );
  XNOR2X1 U4 ( .A(A), .B(B), .Y(n1) );
endmodule


module dff_127 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_126 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_125 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_124 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_123 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_122 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_121 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_120 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_119 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_118 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_117 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_116 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_115 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_114 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_113 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_112 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_111 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_110 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_109 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_108 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_107 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_106 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_105 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_104 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_103 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_102 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_101 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_100 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_99 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_98 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_97 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_96 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_95 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_94 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_93 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_92 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_91 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_90 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_89 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_88 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_87 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_86 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_85 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_84 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_83 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_82 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_81 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_80 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_79 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_78 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_77 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_76 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_75 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_74 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_73 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_72 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_71 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_70 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_69 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_68 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_67 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_66 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_65 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_64 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_63 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_62 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_61 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_60 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_59 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_58 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_57 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_56 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_55 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_54 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_53 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_52 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_51 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_50 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_49 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_48 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_47 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_46 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_45 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_44 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_43 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_42 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_41 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_40 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_39 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_38 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_37 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_36 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_35 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_34 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_33 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_32 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_31 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_30 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_29 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_28 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_27 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_26 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_25 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_24 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_23 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_22 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_21 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_20 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_19 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_18 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_17 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_16 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_15 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_14 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_13 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_12 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_11 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_10 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_9 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_8 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_7 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_6 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_5 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_4 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_3 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_2 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_1 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_0 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module pfa_15 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n4, n2, n3;

  INVX1 U1 ( .A(Cin), .Y(n3) );
  INVX1 U2 ( .A(n2), .Y(P) );
  INVX1 U3 ( .A(n2), .Y(n4) );
  AND2X2 U4 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U5 ( .A(A), .B(B), .Y(n2) );
  XNOR2X1 U6 ( .A(n4), .B(n3), .Y(S) );
endmodule


module pfa_14 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n2;

  XOR2X1 U1 ( .A(B), .B(A), .Y(P) );
  BUFX2 U2 ( .A(P), .Y(n2) );
  AND2X2 U3 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U4 ( .A(Cin), .B(n2), .Y(S) );
endmodule


module pfa_13 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n2, n3, n4;

  XNOR2X1 U1 ( .A(n1), .B(A), .Y(P) );
  INVX1 U2 ( .A(B), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(n2) );
  BUFX2 U4 ( .A(A), .Y(n3) );
  AND2X2 U5 ( .A(B), .B(A), .Y(G) );
  XOR2X1 U6 ( .A(n3), .B(n2), .Y(n4) );
  XOR2X1 U7 ( .A(Cin), .B(n4), .Y(S) );
endmodule


module pfa_12 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n4, n1, n3;

  INVX1 U1 ( .A(P), .Y(n1) );
  INVX1 U2 ( .A(n3), .Y(P) );
  INVX1 U3 ( .A(n1), .Y(n4) );
  XNOR2X1 U4 ( .A(A), .B(B), .Y(n3) );
  AND2X2 U5 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U6 ( .A(Cin), .B(n4), .Y(S) );
endmodule


module pfa_11 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n3;

  INVX1 U1 ( .A(n3), .Y(n1) );
  XOR2X1 U2 ( .A(Cin), .B(n1), .Y(S) );
  XOR2X1 U3 ( .A(B), .B(A), .Y(P) );
  INVX1 U4 ( .A(P), .Y(n3) );
  AND2X2 U5 ( .A(B), .B(A), .Y(G) );
endmodule


module pfa_10 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n2, n3;

  INVX2 U1 ( .A(A), .Y(n2) );
  XNOR2X1 U2 ( .A(B), .B(n2), .Y(P) );
  BUFX2 U3 ( .A(P), .Y(n3) );
  AND2X2 U4 ( .A(B), .B(A), .Y(G) );
  XOR2X1 U5 ( .A(Cin), .B(n3), .Y(S) );
endmodule


module pfa_9 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n2;

  XOR2X1 U1 ( .A(A), .B(B), .Y(P) );
  BUFX2 U2 ( .A(P), .Y(n2) );
  AND2X2 U3 ( .A(B), .B(A), .Y(G) );
  XOR2X1 U4 ( .A(Cin), .B(n2), .Y(S) );
endmodule


module pfa_8 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n3;

  BUFX2 U1 ( .A(P), .Y(n1) );
  XOR2X1 U2 ( .A(B), .B(A), .Y(P) );
  INVX1 U3 ( .A(n1), .Y(n3) );
  XNOR2X1 U4 ( .A(Cin), .B(n3), .Y(S) );
  AND2X2 U5 ( .A(A), .B(B), .Y(G) );
endmodule


module pfa_7 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n2;

  XOR2X1 U1 ( .A(B), .B(A), .Y(P) );
  BUFX2 U2 ( .A(P), .Y(n2) );
  XOR2X1 U3 ( .A(Cin), .B(n2), .Y(S) );
  AND2X2 U4 ( .A(A), .B(B), .Y(G) );
endmodule


module pfa_6 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n2, n4, n5;

  INVX1 U1 ( .A(B), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(n2) );
  XOR2X1 U3 ( .A(n2), .B(A), .Y(P) );
  XOR2X1 U4 ( .A(Cin), .B(n4), .Y(S) );
  INVX1 U5 ( .A(n5), .Y(n4) );
  INVX1 U6 ( .A(P), .Y(n5) );
  AND2X2 U7 ( .A(A), .B(B), .Y(G) );
endmodule


module pfa_5 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n2, n3, n4, n5;

  INVX1 U1 ( .A(n4), .Y(n3) );
  INVX2 U2 ( .A(n5), .Y(P) );
  INVX1 U3 ( .A(B), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n2) );
  XOR2X1 U5 ( .A(Cin), .B(n3), .Y(S) );
  AND2X2 U6 ( .A(A), .B(B), .Y(G) );
  INVX1 U7 ( .A(P), .Y(n4) );
  XNOR2X1 U8 ( .A(n2), .B(A), .Y(n5) );
endmodule


module pfa_4 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n2, n3, n4, n5;

  XOR2X1 U1 ( .A(n2), .B(n5), .Y(P) );
  BUFX2 U2 ( .A(A), .Y(n2) );
  BUFX2 U3 ( .A(P), .Y(n3) );
  INVX1 U4 ( .A(B), .Y(n4) );
  INVX1 U5 ( .A(n4), .Y(n5) );
  AND2X2 U6 ( .A(B), .B(A), .Y(G) );
  XOR2X1 U7 ( .A(Cin), .B(n3), .Y(S) );
endmodule


module pfa_3 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U1 ( .A(A), .B(B), .Y(P) );
  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  AND2X2 U3 ( .A(A), .B(B), .Y(G) );
endmodule


module pfa_2 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  XNOR2X1 U1 ( .A(Cin), .B(n1), .Y(S) );
  INVX1 U2 ( .A(n1), .Y(P) );
  AND2X2 U3 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U4 ( .A(A), .B(B), .Y(n1) );
endmodule


module pfa_1 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n2;

  INVX1 U1 ( .A(A), .Y(n1) );
  XNOR2X1 U2 ( .A(B), .B(n1), .Y(P) );
  BUFX2 U3 ( .A(P), .Y(n2) );
  AND2X2 U4 ( .A(B), .B(A), .Y(G) );
  XOR2X1 U5 ( .A(Cin), .B(n2), .Y(S) );
endmodule


module pfa_0 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U2 ( .A(Cin), .B(n1), .Y(S) );
  XNOR2X1 U3 ( .A(A), .B(B), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(P) );
endmodule


module dff_159 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_158 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_157 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_156 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_155 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_154 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_153 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_152 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_151 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_150 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_149 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_148 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_147 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_146 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_145 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_144 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_143 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_142 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_141 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_140 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_139 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_138 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_137 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_136 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_135 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_134 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_133 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_132 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_131 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_130 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_129 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_128 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module CLA4_23 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, Cout, P, G, .S({\S<3> , \S<2> , \S<1> , \S<0> }
        ) );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output Cout, P, G, \S<3> , \S<2> , \S<1> , \S<0> ;
  wire   p0, g0, p1, g1, p2, g2, c3, p3, g3, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n13, n14, n15, n16, n17, n18, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29;

  pfa_95 bit0 ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(p0), .G(g0)
         );
  pfa_94 bit1 ( .A(\A<1> ), .B(\B<1> ), .Cin(n17), .S(\S<1> ), .P(p1), .G(g1)
         );
  pfa_93 bit2 ( .A(\A<2> ), .B(\B<2> ), .Cin(n14), .S(\S<2> ), .P(p2), .G(g2)
         );
  pfa_92 bit3 ( .A(\A<3> ), .B(\B<3> ), .Cin(c3), .S(\S<3> ), .P(p3), .G(g3)
         );
  INVX1 U1 ( .A(p2), .Y(n22) );
  INVX1 U2 ( .A(g3), .Y(n24) );
  INVX1 U3 ( .A(Cin), .Y(n28) );
  INVX1 U4 ( .A(g2), .Y(n21) );
  OR2X2 U5 ( .A(p2), .B(g2), .Y(n1) );
  AND2X2 U6 ( .A(Cin), .B(p0), .Y(n2) );
  INVX1 U7 ( .A(n2), .Y(n3) );
  OR2X2 U8 ( .A(g1), .B(g2), .Y(n4) );
  INVX1 U9 ( .A(n4), .Y(n5) );
  BUFX2 U10 ( .A(n23), .Y(n6) );
  AND2X2 U11 ( .A(p1), .B(g0), .Y(n7) );
  INVX1 U12 ( .A(n7), .Y(n8) );
  AND2X2 U13 ( .A(n5), .B(n8), .Y(n9) );
  INVX1 U14 ( .A(n9), .Y(n10) );
  AND2X2 U15 ( .A(n24), .B(n6), .Y(n11) );
  INVX1 U16 ( .A(n11), .Y(G) );
  INVX1 U17 ( .A(n11), .Y(n13) );
  INVX1 U18 ( .A(n18), .Y(n14) );
  INVX1 U19 ( .A(n14), .Y(n15) );
  AND2X2 U20 ( .A(n3), .B(n20), .Y(n16) );
  INVX1 U21 ( .A(n16), .Y(n17) );
  AOI21X1 U22 ( .A(n17), .B(p1), .C(g1), .Y(n18) );
  INVX1 U23 ( .A(n13), .Y(n27) );
  AND2X2 U24 ( .A(n26), .B(n25), .Y(P) );
  INVX1 U25 ( .A(P), .Y(n29) );
  AND2X1 U26 ( .A(p3), .B(p2), .Y(n25) );
  INVX2 U27 ( .A(g0), .Y(n20) );
  OAI21X1 U28 ( .A(n15), .B(n22), .C(n21), .Y(c3) );
  NAND3X1 U29 ( .A(n10), .B(n1), .C(p3), .Y(n23) );
  AND2X2 U30 ( .A(p1), .B(p0), .Y(n26) );
  OAI21X1 U31 ( .A(n29), .B(n28), .C(n27), .Y(Cout) );
endmodule


module CLA4_22 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, Cout, P, G, .S({\S<3> , \S<2> , \S<1> , \S<0> }
        ) );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output Cout, P, G, \S<3> , \S<2> , \S<1> , \S<0> ;
  wire   p0, g0, p1, g1, p2, g2, p3, g3, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35;

  pfa_91 bit0 ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(p0), .G(g0)
         );
  pfa_90 bit1 ( .A(\A<1> ), .B(\B<1> ), .Cin(n27), .S(\S<1> ), .P(p1), .G(g1)
         );
  pfa_89 bit2 ( .A(\A<2> ), .B(\B<2> ), .Cin(n5), .S(\S<2> ), .P(p2), .G(g2)
         );
  pfa_88 bit3 ( .A(\A<3> ), .B(\B<3> ), .Cin(n3), .S(\S<3> ), .P(p3), .G(g3)
         );
  INVX1 U1 ( .A(g0), .Y(n28) );
  INVX1 U2 ( .A(g1), .Y(n30) );
  INVX1 U3 ( .A(g2), .Y(n31) );
  INVX1 U4 ( .A(g3), .Y(n35) );
  INVX1 U5 ( .A(n22), .Y(G) );
  AND2X2 U6 ( .A(p1), .B(p0), .Y(n19) );
  AND2X2 U7 ( .A(n31), .B(n29), .Y(n2) );
  INVX1 U8 ( .A(n2), .Y(n3) );
  AND2X2 U9 ( .A(n30), .B(n12), .Y(n4) );
  INVX1 U10 ( .A(n4), .Y(n5) );
  AND2X2 U11 ( .A(n28), .B(n10), .Y(n6) );
  AND2X2 U12 ( .A(p3), .B(n34), .Y(n7) );
  INVX1 U13 ( .A(n7), .Y(n8) );
  AND2X2 U14 ( .A(Cin), .B(p0), .Y(n9) );
  INVX1 U15 ( .A(n9), .Y(n10) );
  AND2X2 U16 ( .A(p1), .B(n26), .Y(n11) );
  INVX1 U17 ( .A(n11), .Y(n12) );
  INVX1 U18 ( .A(n33), .Y(n13) );
  INVX1 U19 ( .A(n13), .Y(n14) );
  AND2X1 U20 ( .A(Cin), .B(P), .Y(n15) );
  INVX1 U21 ( .A(n15), .Y(n16) );
  AND2X1 U22 ( .A(p3), .B(p2), .Y(n17) );
  INVX1 U23 ( .A(n17), .Y(n18) );
  INVX1 U24 ( .A(n19), .Y(n20) );
  INVX1 U25 ( .A(n23), .Y(n21) );
  AND2X2 U26 ( .A(n8), .B(n35), .Y(n22) );
  INVX1 U27 ( .A(n22), .Y(n23) );
  OR2X2 U28 ( .A(n18), .B(n20), .Y(n24) );
  INVX1 U29 ( .A(n24), .Y(P) );
  INVX1 U30 ( .A(n6), .Y(n26) );
  INVX1 U31 ( .A(n6), .Y(n27) );
  INVX1 U32 ( .A(p2), .Y(n32) );
  OAI21X1 U33 ( .A(g1), .B(n11), .C(p2), .Y(n29) );
  AOI21X1 U34 ( .A(p1), .B(g0), .C(g1), .Y(n33) );
  OAI21X1 U35 ( .A(n14), .B(n32), .C(n31), .Y(n34) );
  NAND2X1 U36 ( .A(n21), .B(n16), .Y(Cout) );
endmodule


module CLA4_21 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, Cout, P, G, .S({\S<3> , \S<2> , \S<1> , \S<0> }
        ) );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output Cout, P, G, \S<3> , \S<2> , \S<1> , \S<0> ;
  wire   n39, p0, g0, p1, g1, p2, g2, p3, g3, n1, n3, n4, n5, n6, n8, n9, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35;

  pfa_87 bit0 ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(p0), .G(g0)
         );
  pfa_86 bit1 ( .A(\A<1> ), .B(\B<1> ), .Cin(n21), .S(n39), .P(p1), .G(g1) );
  pfa_85 bit2 ( .A(\A<2> ), .B(\B<2> ), .Cin(n22), .S(\S<2> ), .P(p2), .G(g2)
         );
  pfa_84 bit3 ( .A(\A<3> ), .B(\B<3> ), .Cin(n19), .S(\S<3> ), .P(p3), .G(g3)
         );
  AOI21X1 U12 ( .A(Cin), .B(P), .C(G), .Y(n34) );
  AOI21X1 U13 ( .A(p3), .B(n32), .C(g3), .Y(n33) );
  OAI21X1 U14 ( .A(n17), .B(n35), .C(n27), .Y(n32) );
  AOI21X1 U15 ( .A(g0), .B(p1), .C(g1), .Y(n31) );
  NAND3X1 U16 ( .A(p3), .B(p2), .C(n29), .Y(n30) );
  INVX1 U1 ( .A(g2), .Y(n27) );
  AND2X1 U2 ( .A(Cin), .B(p0), .Y(n5) );
  INVX1 U3 ( .A(p1), .Y(n25) );
  INVX1 U4 ( .A(g1), .Y(n24) );
  INVX1 U5 ( .A(p2), .Y(n35) );
  INVX2 U6 ( .A(n39), .Y(n1) );
  INVX4 U7 ( .A(n1), .Y(\S<1> ) );
  INVX1 U8 ( .A(n21), .Y(n26) );
  AND2X2 U9 ( .A(p2), .B(n28), .Y(n3) );
  INVX1 U10 ( .A(n3), .Y(n4) );
  INVX1 U11 ( .A(n5), .Y(n6) );
  AND2X1 U17 ( .A(p1), .B(p0), .Y(n29) );
  BUFX2 U18 ( .A(n30), .Y(n8) );
  INVX1 U19 ( .A(n8), .Y(P) );
  BUFX2 U20 ( .A(n33), .Y(n9) );
  INVX1 U21 ( .A(n9), .Y(G) );
  BUFX2 U22 ( .A(n34), .Y(n16) );
  INVX1 U23 ( .A(n16), .Y(Cout) );
  BUFX2 U24 ( .A(n31), .Y(n17) );
  AND2X2 U25 ( .A(n27), .B(n4), .Y(n18) );
  INVX1 U26 ( .A(n18), .Y(n19) );
  AND2X2 U27 ( .A(n6), .B(n23), .Y(n20) );
  INVX1 U28 ( .A(n20), .Y(n21) );
  OAI21X1 U29 ( .A(n26), .B(n25), .C(n24), .Y(n22) );
  INVX2 U30 ( .A(g0), .Y(n23) );
  OAI21X1 U31 ( .A(n26), .B(n25), .C(n24), .Y(n28) );
endmodule


module CLA4_20 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, Cout, P, G, .S({\S<3> , \S<2> , \S<1> , \S<0> }
        ) );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output Cout, P, G, \S<3> , \S<2> , \S<1> , \S<0> ;
  wire   p0, g0, p1, g1, p2, g2, c3, p3, g3, n1, n2, n3, n4, n5, n8, n9, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29;

  pfa_83 bit0 ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(p0), .G(g0)
         );
  pfa_82 bit1 ( .A(\A<1> ), .B(\B<1> ), .Cin(n9), .S(\S<1> ), .P(p1), .G(g1)
         );
  pfa_81 bit2 ( .A(\A<2> ), .B(\B<2> ), .Cin(n21), .S(\S<2> ), .P(p2), .G(g2)
         );
  pfa_80 bit3 ( .A(\A<3> ), .B(\B<3> ), .Cin(c3), .S(\S<3> ), .P(p3), .G(g3)
         );
  AOI21X1 U12 ( .A(Cin), .B(P), .C(G), .Y(n27) );
  AOI21X1 U13 ( .A(p3), .B(n25), .C(g3), .Y(n26) );
  OAI21X1 U14 ( .A(n8), .B(n28), .C(n29), .Y(n25) );
  AOI21X1 U15 ( .A(g0), .B(p1), .C(g1), .Y(n24) );
  NAND3X1 U16 ( .A(p3), .B(p2), .C(n22), .Y(n23) );
  INVX1 U1 ( .A(g0), .Y(n17) );
  INVX1 U2 ( .A(p2), .Y(n28) );
  INVX1 U3 ( .A(g2), .Y(n29) );
  INVX1 U4 ( .A(g1), .Y(n18) );
  INVX1 U5 ( .A(p1), .Y(n19) );
  AND2X1 U6 ( .A(p1), .B(p0), .Y(n22) );
  AND2X1 U7 ( .A(p0), .B(Cin), .Y(n1) );
  INVX1 U8 ( .A(n1), .Y(n2) );
  BUFX2 U9 ( .A(n23), .Y(n3) );
  INVX1 U10 ( .A(n3), .Y(P) );
  BUFX2 U11 ( .A(n26), .Y(n4) );
  INVX1 U17 ( .A(n4), .Y(G) );
  BUFX2 U18 ( .A(n27), .Y(n5) );
  INVX1 U19 ( .A(n5), .Y(Cout) );
  BUFX2 U20 ( .A(n24), .Y(n8) );
  INVX1 U21 ( .A(n16), .Y(n9) );
  AND2X2 U22 ( .A(n17), .B(n2), .Y(n16) );
  OAI21X1 U23 ( .A(n16), .B(n19), .C(n18), .Y(n21) );
  INVX2 U24 ( .A(n21), .Y(n20) );
  OAI21X1 U25 ( .A(n20), .B(n28), .C(n29), .Y(c3) );
endmodule


module CLA4_19 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, Cout, P, G, .S({\S<3> , \S<2> , \S<1> , \S<0> }
        ) );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output Cout, P, G, \S<3> , \S<2> , \S<1> , \S<0> ;
  wire   p0, g0, p1, g1, p2, g2, c3, p3, g3, n1, n2, n4, n5, n6, n7, n8, n9,
         n10, n11, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n28;

  pfa_79 bit0 ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(p0), .G(g0)
         );
  pfa_78 bit1 ( .A(\A<1> ), .B(\B<1> ), .Cin(n5), .S(\S<1> ), .P(p1), .G(g1)
         );
  pfa_77 bit2 ( .A(\A<2> ), .B(\B<2> ), .Cin(n28), .S(\S<2> ), .P(p2), .G(g2)
         );
  pfa_76 bit3 ( .A(\A<3> ), .B(\B<3> ), .Cin(c3), .S(\S<3> ), .P(p3), .G(g3)
         );
  INVX1 U1 ( .A(g0), .Y(n15) );
  INVX1 U2 ( .A(p2), .Y(n20) );
  INVX1 U3 ( .A(g2), .Y(n19) );
  INVX1 U4 ( .A(Cin), .Y(n26) );
  BUFX2 U5 ( .A(p1), .Y(n1) );
  INVX1 U6 ( .A(g1), .Y(n16) );
  AND2X2 U7 ( .A(n23), .B(n8), .Y(n2) );
  INVX1 U8 ( .A(n2), .Y(G) );
  AND2X2 U9 ( .A(n15), .B(n7), .Y(n4) );
  INVX1 U10 ( .A(n4), .Y(n5) );
  AND2X2 U11 ( .A(Cin), .B(p0), .Y(n6) );
  INVX1 U12 ( .A(n6), .Y(n7) );
  INVX1 U13 ( .A(n10), .Y(n8) );
  AND2X2 U14 ( .A(n22), .B(p3), .Y(n10) );
  BUFX2 U15 ( .A(n21), .Y(n9) );
  INVX1 U16 ( .A(n10), .Y(n11) );
  AND2X2 U17 ( .A(n25), .B(n24), .Y(P) );
  INVX1 U18 ( .A(P), .Y(n13) );
  AND2X2 U19 ( .A(n11), .B(n23), .Y(n14) );
  INVX1 U20 ( .A(g3), .Y(n23) );
  INVX1 U21 ( .A(n1), .Y(n17) );
  OAI21X1 U22 ( .A(n4), .B(n17), .C(n16), .Y(n28) );
  INVX2 U23 ( .A(n28), .Y(n18) );
  OAI21X1 U24 ( .A(n18), .B(n20), .C(n19), .Y(c3) );
  AOI21X1 U25 ( .A(p1), .B(g0), .C(g1), .Y(n21) );
  OAI21X1 U26 ( .A(n9), .B(n20), .C(n19), .Y(n22) );
  AND2X2 U27 ( .A(n1), .B(p0), .Y(n25) );
  AND2X2 U28 ( .A(p3), .B(p2), .Y(n24) );
  OAI21X1 U29 ( .A(n13), .B(n26), .C(n14), .Y(Cout) );
endmodule


module CLA4_18 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, Cout, P, G, .S({\S<3> , \S<2> , \S<1> , \S<0> }
        ) );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output Cout, P, G, \S<3> , \S<2> , \S<1> , \S<0> ;
  wire   p0, g0, p1, g1, p2, g2, c3, p3, g3, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n23,
         n25, n26, n27, n28, n29, n30, n31, n32;

  pfa_75 bit0 ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(p0), .G(g0)
         );
  pfa_74 bit1 ( .A(\A<1> ), .B(\B<1> ), .Cin(n19), .S(\S<1> ), .P(p1), .G(g1)
         );
  pfa_73 bit2 ( .A(\A<2> ), .B(\B<2> ), .Cin(n2), .S(\S<2> ), .P(p2), .G(g2)
         );
  pfa_72 bit3 ( .A(\A<3> ), .B(\B<3> ), .Cin(c3), .S(\S<3> ), .P(p3), .G(g3)
         );
  INVX1 U1 ( .A(g0), .Y(n27) );
  INVX1 U2 ( .A(p2), .Y(n29) );
  INVX1 U3 ( .A(g2), .Y(n28) );
  INVX1 U4 ( .A(g3), .Y(n32) );
  AND2X2 U5 ( .A(Cin), .B(P), .Y(n10) );
  AND2X2 U6 ( .A(n26), .B(n20), .Y(n1) );
  INVX1 U7 ( .A(n1), .Y(n2) );
  AND2X2 U8 ( .A(n27), .B(n5), .Y(n3) );
  AND2X2 U9 ( .A(Cin), .B(p0), .Y(n4) );
  INVX1 U10 ( .A(n4), .Y(n5) );
  AND2X2 U11 ( .A(p1), .B(n18), .Y(n6) );
  INVX1 U12 ( .A(n6), .Y(n7) );
  AND2X1 U13 ( .A(p3), .B(n31), .Y(n8) );
  INVX1 U14 ( .A(n8), .Y(n9) );
  INVX1 U15 ( .A(n10), .Y(n11) );
  AND2X1 U16 ( .A(p3), .B(p2), .Y(n12) );
  INVX1 U17 ( .A(n12), .Y(n13) );
  AND2X1 U18 ( .A(p1), .B(p0), .Y(n14) );
  INVX1 U19 ( .A(n14), .Y(n15) );
  INVX1 U20 ( .A(n30), .Y(n16) );
  INVX1 U21 ( .A(n16), .Y(n17) );
  INVX1 U22 ( .A(n3), .Y(n18) );
  INVX1 U23 ( .A(n3), .Y(n19) );
  INVX1 U24 ( .A(n6), .Y(n20) );
  OR2X2 U25 ( .A(n13), .B(n15), .Y(n21) );
  INVX1 U26 ( .A(n21), .Y(P) );
  AND2X2 U27 ( .A(n32), .B(n9), .Y(n23) );
  INVX1 U28 ( .A(n23), .Y(G) );
  AND2X2 U29 ( .A(n7), .B(n26), .Y(n25) );
  INVX1 U30 ( .A(g1), .Y(n26) );
  OAI21X1 U31 ( .A(n25), .B(n29), .C(n28), .Y(c3) );
  AOI21X1 U32 ( .A(p1), .B(g0), .C(g1), .Y(n30) );
  OAI21X1 U33 ( .A(n17), .B(n29), .C(n28), .Y(n31) );
  NAND2X1 U34 ( .A(n23), .B(n11), .Y(Cout) );
endmodule


module CLA4_17 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, Cout, P, G, .S({\S<3> , \S<2> , \S<1> , \S<0> }
        ) );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output Cout, P, G, \S<3> , \S<2> , \S<1> , \S<0> ;
  wire   p0, g0, p1, g1, p2, g2, p3, g3, n1, n2, n3, n4, n5, n6, n8, n9, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33;

  pfa_71 bit0 ( .A(\A<0> ), .B(\B<0> ), .Cin(n2), .S(\S<0> ), .P(p0), .G(g0)
         );
  pfa_70 bit1 ( .A(\A<1> ), .B(\B<1> ), .Cin(n21), .S(\S<1> ), .P(p1), .G(g1)
         );
  pfa_69 bit2 ( .A(\A<2> ), .B(\B<2> ), .Cin(n1), .S(\S<2> ), .P(p2), .G(g2)
         );
  pfa_68 bit3 ( .A(\A<3> ), .B(\B<3> ), .Cin(n4), .S(\S<3> ), .P(p3), .G(g3)
         );
  AOI21X1 U12 ( .A(n2), .B(P), .C(G), .Y(n32) );
  AOI21X1 U13 ( .A(p3), .B(n30), .C(g3), .Y(n31) );
  OAI21X1 U14 ( .A(n19), .B(n33), .C(n25), .Y(n30) );
  AOI21X1 U15 ( .A(g0), .B(p1), .C(g1), .Y(n29) );
  NAND3X1 U16 ( .A(p3), .B(p2), .C(n27), .Y(n28) );
  INVX1 U1 ( .A(g2), .Y(n25) );
  INVX1 U2 ( .A(g1), .Y(n23) );
  INVX1 U3 ( .A(g0), .Y(n22) );
  INVX1 U4 ( .A(p2), .Y(n33) );
  OAI21X1 U5 ( .A(n24), .B(n20), .C(n23), .Y(n1) );
  BUFX2 U6 ( .A(Cin), .Y(n2) );
  AND2X1 U7 ( .A(Cin), .B(p0), .Y(n5) );
  AND2X2 U8 ( .A(n25), .B(n9), .Y(n3) );
  INVX1 U9 ( .A(n3), .Y(n4) );
  INVX1 U10 ( .A(n5), .Y(n6) );
  AND2X2 U11 ( .A(p2), .B(n26), .Y(n8) );
  INVX1 U17 ( .A(n8), .Y(n9) );
  AND2X1 U18 ( .A(p1), .B(p0), .Y(n27) );
  BUFX2 U19 ( .A(n28), .Y(n16) );
  INVX1 U20 ( .A(n16), .Y(P) );
  BUFX2 U21 ( .A(n31), .Y(n17) );
  INVX1 U22 ( .A(n17), .Y(G) );
  BUFX2 U23 ( .A(n32), .Y(n18) );
  INVX1 U24 ( .A(n18), .Y(Cout) );
  BUFX2 U25 ( .A(n29), .Y(n19) );
  AND2X2 U26 ( .A(n6), .B(n22), .Y(n20) );
  INVX1 U27 ( .A(n20), .Y(n21) );
  INVX2 U28 ( .A(p1), .Y(n24) );
  OAI21X1 U29 ( .A(n24), .B(n20), .C(n23), .Y(n26) );
endmodule


module CLA4_16 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, Cout, P, G, .S({\S<3> , \S<2> , \S<1> , \S<0> }
        ) );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output Cout, P, G, \S<3> , \S<2> , \S<1> , \S<0> ;
  wire   p0, g0, p1, g1, p2, g2, c3, p3, g3, n3, n4, n5, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n31, n32;

  pfa_67 bit0 ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(p0), .G(g0)
         );
  pfa_66 bit1 ( .A(\A<1> ), .B(\B<1> ), .Cin(n31), .S(\S<1> ), .P(p1), .G(g1)
         );
  pfa_65 bit2 ( .A(\A<2> ), .B(\B<2> ), .Cin(n32), .S(\S<2> ), .P(p2), .G(g2)
         );
  pfa_64 bit3 ( .A(\A<3> ), .B(\B<3> ), .Cin(c3), .S(\S<3> ), .P(p3), .G(g3)
         );
  OAI21X1 U9 ( .A(n17), .B(n26), .C(n27), .Y(c3) );
  AOI21X1 U10 ( .A(p1), .B(n31), .C(g1), .Y(n25) );
  AOI21X1 U11 ( .A(Cin), .B(p0), .C(g0), .Y(n24) );
  AOI21X1 U12 ( .A(Cin), .B(P), .C(G), .Y(n23) );
  AOI21X1 U13 ( .A(p3), .B(n21), .C(g3), .Y(n22) );
  OAI21X1 U14 ( .A(n16), .B(n26), .C(n27), .Y(n21) );
  AOI21X1 U15 ( .A(g0), .B(p1), .C(g1), .Y(n20) );
  NAND3X1 U16 ( .A(p3), .B(p2), .C(n18), .Y(n19) );
  INVX1 U1 ( .A(p2), .Y(n26) );
  INVX1 U2 ( .A(g2), .Y(n27) );
  INVX1 U3 ( .A(n17), .Y(n32) );
  AND2X1 U4 ( .A(p1), .B(p0), .Y(n18) );
  BUFX2 U5 ( .A(n19), .Y(n3) );
  INVX1 U6 ( .A(n3), .Y(P) );
  BUFX2 U7 ( .A(n22), .Y(n4) );
  INVX1 U8 ( .A(n4), .Y(G) );
  BUFX2 U17 ( .A(n23), .Y(n5) );
  INVX1 U18 ( .A(n5), .Y(Cout) );
  INVX1 U19 ( .A(n24), .Y(n31) );
  BUFX2 U20 ( .A(n20), .Y(n16) );
  BUFX2 U21 ( .A(n25), .Y(n17) );
endmodule


module CLA4_15 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, Cout, P, G, .S({\S<3> , \S<2> , \S<1> , \S<0> }
        ) );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output Cout, P, G, \S<3> , \S<2> , \S<1> , \S<0> ;
  wire   p0, g0, p1, g1, p2, g2, c3, p3, g3, n1, n3, n4, n6, n7, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n23, n24, n26;

  pfa_63 bit0 ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(p0), .G(g0)
         );
  pfa_62 bit1 ( .A(\A<1> ), .B(\B<1> ), .Cin(n26), .S(\S<1> ), .P(p1), .G(g1)
         );
  pfa_61 bit2 ( .A(\A<2> ), .B(\B<2> ), .Cin(n7), .S(\S<2> ), .P(p2), .G(g2)
         );
  pfa_60 bit3 ( .A(\A<3> ), .B(\B<3> ), .Cin(c3), .S(\S<3> ), .P(p3), .G(g3)
         );
  AOI21X1 U10 ( .A(n26), .B(p1), .C(g1), .Y(n24) );
  AOI21X1 U11 ( .A(Cin), .B(p0), .C(g0), .Y(n23) );
  INVX1 U1 ( .A(p2), .Y(n12) );
  INVX1 U2 ( .A(g2), .Y(n11) );
  INVX1 U3 ( .A(g3), .Y(n17) );
  INVX1 U4 ( .A(G), .Y(n19) );
  INVX1 U5 ( .A(Cin), .Y(n20) );
  BUFX2 U6 ( .A(n13), .Y(n1) );
  INVX1 U7 ( .A(n1), .Y(n14) );
  BUFX2 U8 ( .A(n23), .Y(n3) );
  INVX1 U9 ( .A(n3), .Y(n26) );
  AND2X2 U12 ( .A(n17), .B(n16), .Y(n4) );
  INVX1 U13 ( .A(n4), .Y(G) );
  INVX1 U14 ( .A(P), .Y(n6) );
  INVX1 U15 ( .A(n21), .Y(P) );
  INVX1 U16 ( .A(n10), .Y(n7) );
  BUFX2 U17 ( .A(n24), .Y(n10) );
  OAI21X1 U18 ( .A(n10), .B(n12), .C(n11), .Y(c3) );
  AOI21X1 U19 ( .A(g0), .B(p1), .C(g1), .Y(n13) );
  AND2X2 U20 ( .A(p2), .B(n14), .Y(n15) );
  OAI21X1 U21 ( .A(n15), .B(g2), .C(p3), .Y(n16) );
  AND2X2 U22 ( .A(p0), .B(p1), .Y(n18) );
  NAND3X1 U23 ( .A(p2), .B(n18), .C(p3), .Y(n21) );
  OAI21X1 U24 ( .A(n6), .B(n20), .C(n19), .Y(Cout) );
endmodule


module CLA4_14 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, Cout, P, G, .S({\S<3> , \S<2> , \S<1> , \S<0> }
        ) );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output Cout, P, G, \S<3> , \S<2> , \S<1> , \S<0> ;
  wire   p0, g0, p1, g1, p2, g2, c3, p3, g3, n3, n4, n5, n6, n7, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n25, n26, n28;

  pfa_59 bit0 ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(p0), .G(g0)
         );
  pfa_58 bit1 ( .A(\A<1> ), .B(\B<1> ), .Cin(n28), .S(\S<1> ), .P(p1), .G(g1)
         );
  pfa_57 bit2 ( .A(\A<2> ), .B(\B<2> ), .Cin(n12), .S(\S<2> ), .P(p2), .G(g2)
         );
  pfa_56 bit3 ( .A(\A<3> ), .B(\B<3> ), .Cin(c3), .S(\S<3> ), .P(p3), .G(g3)
         );
  AOI21X1 U10 ( .A(n28), .B(p1), .C(g1), .Y(n26) );
  AOI21X1 U11 ( .A(Cin), .B(p0), .C(g0), .Y(n25) );
  INVX1 U1 ( .A(g2), .Y(n15) );
  INVX1 U2 ( .A(g1), .Y(n17) );
  INVX1 U3 ( .A(g3), .Y(n20) );
  INVX1 U4 ( .A(n5), .Y(G) );
  INVX1 U5 ( .A(p2), .Y(n16) );
  AND2X2 U6 ( .A(g0), .B(p1), .Y(n3) );
  INVX1 U7 ( .A(n3), .Y(n4) );
  AND2X2 U8 ( .A(n20), .B(n19), .Y(n5) );
  AND2X2 U9 ( .A(n17), .B(n4), .Y(n6) );
  INVX1 U12 ( .A(n6), .Y(n7) );
  INVX1 U13 ( .A(Cin), .Y(n22) );
  BUFX2 U14 ( .A(n25), .Y(n10) );
  INVX1 U15 ( .A(n10), .Y(n28) );
  INVX1 U16 ( .A(P), .Y(n11) );
  INVX1 U17 ( .A(n23), .Y(P) );
  INVX1 U18 ( .A(n13), .Y(n12) );
  BUFX2 U19 ( .A(n26), .Y(n13) );
  INVX1 U20 ( .A(G), .Y(n14) );
  OAI21X1 U21 ( .A(n13), .B(n16), .C(n15), .Y(c3) );
  AND2X2 U22 ( .A(p2), .B(n7), .Y(n18) );
  OAI21X1 U23 ( .A(n18), .B(g2), .C(p3), .Y(n19) );
  AND2X2 U24 ( .A(p0), .B(p1), .Y(n21) );
  NAND3X1 U25 ( .A(p2), .B(n21), .C(p3), .Y(n23) );
  OAI21X1 U26 ( .A(n11), .B(n22), .C(n14), .Y(Cout) );
endmodule


module CLA4_13 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, Cout, P, G, .S({\S<3> , \S<2> , \S<1> , \S<0> }
        ) );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output Cout, P, G, \S<3> , \S<2> , \S<1> , \S<0> ;
  wire   p0, g0, p1, g1, p2, g2, p3, g3, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n38;

  pfa_55 bit0 ( .A(\A<0> ), .B(\B<0> ), .Cin(n27), .S(\S<0> ), .P(p0), .G(g0)
         );
  pfa_54 bit1 ( .A(\A<1> ), .B(\B<1> ), .Cin(n6), .S(\S<1> ), .P(p1), .G(g1)
         );
  pfa_53 bit2 ( .A(\A<2> ), .B(\B<2> ), .Cin(n25), .S(\S<2> ), .P(p2), .G(g2)
         );
  pfa_52 bit3 ( .A(\A<3> ), .B(\B<3> ), .Cin(n18), .S(\S<3> ), .P(p3), .G(g3)
         );
  AND2X1 U1 ( .A(n38), .B(p2), .Y(n9) );
  INVX1 U2 ( .A(g2), .Y(n30) );
  AND2X1 U3 ( .A(p1), .B(g0), .Y(n13) );
  INVX1 U4 ( .A(g1), .Y(n31) );
  INVX1 U5 ( .A(g3), .Y(n34) );
  BUFX2 U6 ( .A(p1), .Y(n1) );
  OR2X2 U7 ( .A(n17), .B(n3), .Y(n12) );
  INVX1 U8 ( .A(n1), .Y(n29) );
  INVX1 U9 ( .A(G), .Y(n36) );
  AND2X2 U10 ( .A(n21), .B(n28), .Y(n2) );
  INVX1 U11 ( .A(p3), .Y(n3) );
  INVX1 U12 ( .A(n3), .Y(n4) );
  AND2X2 U13 ( .A(n27), .B(P), .Y(n15) );
  AND2X2 U14 ( .A(n34), .B(n33), .Y(n11) );
  AND2X2 U15 ( .A(n28), .B(n21), .Y(n5) );
  INVX1 U16 ( .A(n5), .Y(n6) );
  AND2X2 U17 ( .A(n31), .B(n14), .Y(n7) );
  INVX1 U18 ( .A(n7), .Y(n8) );
  INVX1 U19 ( .A(n9), .Y(n10) );
  INVX1 U20 ( .A(n13), .Y(n14) );
  INVX1 U21 ( .A(n15), .Y(n16) );
  BUFX2 U22 ( .A(n35), .Y(n17) );
  INVX1 U23 ( .A(n19), .Y(n18) );
  AND2X2 U24 ( .A(n30), .B(n10), .Y(n19) );
  AND2X2 U25 ( .A(Cin), .B(p0), .Y(n20) );
  INVX1 U26 ( .A(n20), .Y(n21) );
  INVX1 U27 ( .A(n12), .Y(P) );
  INVX1 U28 ( .A(n11), .Y(G) );
  AND2X2 U29 ( .A(n21), .B(n28), .Y(n24) );
  INVX1 U30 ( .A(g0), .Y(n28) );
  OAI21X1 U31 ( .A(n2), .B(n29), .C(n31), .Y(n25) );
  INVX1 U32 ( .A(Cin), .Y(n26) );
  INVX1 U33 ( .A(n26), .Y(n27) );
  OAI21X1 U34 ( .A(n24), .B(n29), .C(n31), .Y(n38) );
  AND2X2 U35 ( .A(p2), .B(n8), .Y(n32) );
  OAI21X1 U36 ( .A(n32), .B(g2), .C(n4), .Y(n33) );
  NAND3X1 U37 ( .A(n1), .B(p0), .C(p2), .Y(n35) );
  NAND2X1 U38 ( .A(n36), .B(n16), .Y(Cout) );
endmodule


module CLA4_12 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, Cout, P, G, .S({\S<3> , \S<2> , \S<1> , \S<0> }
        ) );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output Cout, P, G, \S<3> , \S<2> , \S<1> , \S<0> ;
  wire   p0, g0, p1, g1, p2, g2, p3, g3, n1, n2, n3, n4, n5, n6, n8, n9, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43;

  pfa_51 bit0 ( .A(\A<0> ), .B(\B<0> ), .Cin(n5), .S(\S<0> ), .P(p0), .G(g0)
         );
  pfa_50 bit1 ( .A(\A<1> ), .B(\B<1> ), .Cin(n31), .S(\S<1> ), .P(p1), .G(g1)
         );
  pfa_49 bit2 ( .A(\A<2> ), .B(\B<2> ), .Cin(n9), .S(\S<2> ), .P(p2), .G(g2)
         );
  pfa_48 bit3 ( .A(\A<3> ), .B(\B<3> ), .Cin(n25), .S(\S<3> ), .P(p3), .G(g3)
         );
  AND2X2 U1 ( .A(p1), .B(p0), .Y(n37) );
  AOI21X1 U12 ( .A(n5), .B(P), .C(G), .Y(n42) );
  AOI21X1 U13 ( .A(p3), .B(n40), .C(g3), .Y(n41) );
  OAI21X1 U14 ( .A(n24), .B(n43), .C(n35), .Y(n40) );
  AOI21X1 U15 ( .A(g0), .B(p1), .C(g1), .Y(n39) );
  NAND3X1 U16 ( .A(p3), .B(n1), .C(n37), .Y(n38) );
  INVX1 U2 ( .A(g1), .Y(n34) );
  INVX1 U3 ( .A(g2), .Y(n35) );
  INVX1 U4 ( .A(n1), .Y(n43) );
  INVX1 U5 ( .A(n21), .Y(Cout) );
  BUFX2 U6 ( .A(p2), .Y(n1) );
  OR2X2 U7 ( .A(g0), .B(n29), .Y(n22) );
  AND2X2 U8 ( .A(p2), .B(g1), .Y(n16) );
  BUFX2 U9 ( .A(n26), .Y(n2) );
  INVX1 U10 ( .A(n26), .Y(n3) );
  INVX1 U11 ( .A(Cin), .Y(n4) );
  INVX1 U17 ( .A(n4), .Y(n5) );
  AND2X2 U18 ( .A(Cin), .B(p0), .Y(n26) );
  AND2X2 U19 ( .A(p1), .B(n31), .Y(n6) );
  AND2X2 U20 ( .A(n34), .B(n18), .Y(n8) );
  INVX1 U21 ( .A(n8), .Y(n9) );
  INVX1 U22 ( .A(n16), .Y(n17) );
  INVX1 U23 ( .A(n6), .Y(n18) );
  BUFX2 U24 ( .A(n32), .Y(n19) );
  BUFX2 U25 ( .A(n38), .Y(n20) );
  INVX1 U26 ( .A(n20), .Y(P) );
  BUFX2 U27 ( .A(n42), .Y(n21) );
  INVX1 U28 ( .A(n41), .Y(G) );
  INVX1 U29 ( .A(n22), .Y(n23) );
  BUFX2 U30 ( .A(n39), .Y(n24) );
  BUFX2 U31 ( .A(n36), .Y(n25) );
  INVX1 U32 ( .A(n2), .Y(n27) );
  AND2X2 U33 ( .A(n35), .B(n17), .Y(n28) );
  INVX1 U34 ( .A(n28), .Y(n29) );
  AND2X2 U35 ( .A(n3), .B(n33), .Y(n30) );
  INVX1 U36 ( .A(n30), .Y(n31) );
  AOI21X1 U37 ( .A(p1), .B(n1), .C(n29), .Y(n32) );
  AOI21X1 U38 ( .A(n23), .B(n27), .C(n19), .Y(n36) );
  INVX2 U39 ( .A(g0), .Y(n33) );
endmodule


module CLA4_11 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, Cout, P, G, .S({\S<3> , \S<2> , \S<1> , \S<0> }
        ) );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output Cout, P, G, \S<3> , \S<2> , \S<1> , \S<0> ;
  wire   p0, g0, p1, g1, p2, g2, c3, p3, g3, n1, n3, n4, n6, n7, n10, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n26, n27, n28;

  pfa_47 bit0 ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(p0), .G(g0)
         );
  pfa_46 bit1 ( .A(\A<1> ), .B(\B<1> ), .Cin(n28), .S(\S<1> ), .P(p1), .G(g1)
         );
  pfa_45 bit2 ( .A(\A<2> ), .B(\B<2> ), .Cin(n13), .S(\S<2> ), .P(p2), .G(g2)
         );
  pfa_44 bit3 ( .A(\A<3> ), .B(\B<3> ), .Cin(c3), .S(\S<3> ), .P(p3), .G(g3)
         );
  AOI21X1 U10 ( .A(n28), .B(p1), .C(g1), .Y(n27) );
  AOI21X1 U11 ( .A(Cin), .B(p0), .C(g0), .Y(n26) );
  INVX1 U1 ( .A(g1), .Y(n17) );
  INVX1 U2 ( .A(p2), .Y(n16) );
  INVX1 U3 ( .A(g2), .Y(n15) );
  INVX1 U4 ( .A(g3), .Y(n20) );
  INVX1 U5 ( .A(G), .Y(n22) );
  INVX1 U6 ( .A(Cin), .Y(n23) );
  AND2X2 U7 ( .A(n17), .B(n7), .Y(n1) );
  INVX1 U8 ( .A(n1), .Y(n3) );
  AND2X2 U9 ( .A(n20), .B(n19), .Y(n4) );
  INVX1 U12 ( .A(n4), .Y(G) );
  AND2X1 U13 ( .A(g0), .B(p1), .Y(n6) );
  INVX1 U14 ( .A(n6), .Y(n7) );
  BUFX2 U15 ( .A(n26), .Y(n10) );
  INVX1 U16 ( .A(n10), .Y(n28) );
  INVX1 U17 ( .A(n24), .Y(P) );
  INVX1 U18 ( .A(P), .Y(n12) );
  INVX1 U19 ( .A(n14), .Y(n13) );
  BUFX2 U20 ( .A(n27), .Y(n14) );
  OAI21X1 U21 ( .A(n14), .B(n16), .C(n15), .Y(c3) );
  AND2X2 U22 ( .A(p2), .B(n3), .Y(n18) );
  OAI21X1 U23 ( .A(n18), .B(g2), .C(p3), .Y(n19) );
  AND2X2 U24 ( .A(p0), .B(p1), .Y(n21) );
  NAND3X1 U25 ( .A(p2), .B(n21), .C(p3), .Y(n24) );
  OAI21X1 U26 ( .A(n12), .B(n23), .C(n22), .Y(Cout) );
endmodule


module CLA4_10 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, Cout, P, G, .S({\S<3> , \S<2> , \S<1> , \S<0> }
        ) );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output Cout, P, G, \S<3> , \S<2> , \S<1> , \S<0> ;
  wire   p0, g0, p1, g1, p2, g2, c3, p3, g3, n1, n3, n4, n5, n6, n7, n10, n11,
         n12, n14, n15, n16, n17, n18, n19, n20, n21, n22, n24, n25, n27;

  pfa_43 bit0 ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(p0), .G(g0)
         );
  pfa_42 bit1 ( .A(\A<1> ), .B(\B<1> ), .Cin(n27), .S(\S<1> ), .P(p1), .G(g1)
         );
  pfa_41 bit2 ( .A(\A<2> ), .B(\B<2> ), .Cin(n10), .S(\S<2> ), .P(p2), .G(g2)
         );
  pfa_40 bit3 ( .A(\A<3> ), .B(\B<3> ), .Cin(c3), .S(\S<3> ), .P(p3), .G(g3)
         );
  AOI21X1 U10 ( .A(n27), .B(p1), .C(g1), .Y(n25) );
  AOI21X1 U11 ( .A(Cin), .B(p0), .C(g0), .Y(n24) );
  INVX1 U1 ( .A(g2), .Y(n17) );
  INVX1 U2 ( .A(p2), .Y(n14) );
  AND2X2 U3 ( .A(p3), .B(n5), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  AND2X2 U5 ( .A(n16), .B(n17), .Y(n4) );
  INVX1 U6 ( .A(n4), .Y(n5) );
  INVX1 U7 ( .A(Cin), .Y(n21) );
  BUFX2 U8 ( .A(n24), .Y(n6) );
  INVX1 U9 ( .A(n6), .Y(n27) );
  INVX1 U12 ( .A(P), .Y(n7) );
  INVX1 U13 ( .A(n11), .Y(n10) );
  BUFX2 U14 ( .A(n25), .Y(n11) );
  AND2X2 U15 ( .A(n3), .B(n18), .Y(n12) );
  INVX1 U16 ( .A(n12), .Y(G) );
  INVX1 U17 ( .A(G), .Y(n20) );
  INVX1 U18 ( .A(n22), .Y(P) );
  OAI21X1 U19 ( .A(n11), .B(n14), .C(n17), .Y(c3) );
  INVX2 U20 ( .A(g3), .Y(n18) );
  AND2X2 U21 ( .A(g0), .B(p1), .Y(n15) );
  OAI21X1 U22 ( .A(n15), .B(g1), .C(p2), .Y(n16) );
  AND2X2 U23 ( .A(p2), .B(p1), .Y(n19) );
  NAND3X1 U24 ( .A(p0), .B(p3), .C(n19), .Y(n22) );
  OAI21X1 U25 ( .A(n7), .B(n21), .C(n20), .Y(Cout) );
endmodule


module CLA4_9 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, Cout, P, G, .S({\S<3> , \S<2> , \S<1> , \S<0> }
        ) );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output Cout, P, G, \S<3> , \S<2> , \S<1> , \S<0> ;
  wire   p0, g0, p1, g1, p2, g2, p3, g3, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n11, n12, n13, n14, n15, n16, n17, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n35;

  pfa_39 bit0 ( .A(\A<0> ), .B(\B<0> ), .Cin(n23), .S(\S<0> ), .P(p0), .G(g0)
         );
  pfa_38 bit1 ( .A(\A<1> ), .B(\B<1> ), .Cin(n20), .S(\S<1> ), .P(p1), .G(g1)
         );
  pfa_37 bit2 ( .A(\A<2> ), .B(\B<2> ), .Cin(n21), .S(\S<2> ), .P(p2), .G(g2)
         );
  pfa_36 bit3 ( .A(\A<3> ), .B(\B<3> ), .Cin(n15), .S(\S<3> ), .P(p3), .G(g3)
         );
  INVX1 U1 ( .A(g1), .Y(n27) );
  INVX1 U2 ( .A(g0), .Y(n24) );
  INVX1 U3 ( .A(g3), .Y(n30) );
  BUFX2 U4 ( .A(p1), .Y(n1) );
  AND2X1 U5 ( .A(p1), .B(g0), .Y(n11) );
  AND2X2 U6 ( .A(p3), .B(n32), .Y(P) );
  INVX1 U7 ( .A(n1), .Y(n25) );
  AND2X2 U8 ( .A(n30), .B(n29), .Y(n17) );
  AND2X2 U9 ( .A(p2), .B(n35), .Y(n8) );
  AND2X2 U10 ( .A(n24), .B(n7), .Y(n2) );
  INVX1 U11 ( .A(n2), .Y(n3) );
  AND2X2 U12 ( .A(n27), .B(n12), .Y(n4) );
  INVX1 U13 ( .A(n4), .Y(n5) );
  AND2X2 U14 ( .A(Cin), .B(p0), .Y(n6) );
  INVX1 U15 ( .A(n6), .Y(n7) );
  INVX1 U16 ( .A(n8), .Y(n9) );
  INVX1 U17 ( .A(n11), .Y(n12) );
  AND2X1 U18 ( .A(n23), .B(P), .Y(n13) );
  INVX1 U19 ( .A(n13), .Y(n14) );
  INVX1 U20 ( .A(n16), .Y(n15) );
  AND2X2 U21 ( .A(n9), .B(n26), .Y(n16) );
  INVX1 U22 ( .A(n17), .Y(G) );
  INVX1 U23 ( .A(n3), .Y(n19) );
  INVX1 U24 ( .A(n19), .Y(n20) );
  OAI21X1 U25 ( .A(n19), .B(n25), .C(n27), .Y(n21) );
  INVX1 U26 ( .A(Cin), .Y(n22) );
  INVX1 U27 ( .A(n22), .Y(n23) );
  INVX1 U28 ( .A(G), .Y(n33) );
  OAI21X1 U29 ( .A(n2), .B(n25), .C(n27), .Y(n35) );
  INVX2 U30 ( .A(g2), .Y(n26) );
  AND2X2 U31 ( .A(p2), .B(n5), .Y(n28) );
  OAI21X1 U32 ( .A(n28), .B(g2), .C(p3), .Y(n29) );
  AND2X2 U33 ( .A(n1), .B(p0), .Y(n31) );
  AND2X2 U34 ( .A(p2), .B(n31), .Y(n32) );
  NAND2X1 U35 ( .A(n33), .B(n14), .Y(Cout) );
endmodule


module CLA4_8 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, Cout, P, G, .S({\S<3> , \S<2> , \S<1> , \S<0> }
        ) );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output Cout, P, G, \S<3> , \S<2> , \S<1> , \S<0> ;
  wire   p0, g0, p1, g1, p2, g2, p3, g3, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n11, n12, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n32, n33, n34, n35;

  pfa_35 bit0 ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(p0), .G(g0)
         );
  pfa_34 bit1 ( .A(\A<1> ), .B(\B<1> ), .Cin(n18), .S(\S<1> ), .P(p1), .G(g1)
         );
  pfa_33 bit2 ( .A(\A<2> ), .B(\B<2> ), .Cin(n30), .S(\S<2> ), .P(p2), .G(g2)
         );
  pfa_32 bit3 ( .A(\A<3> ), .B(\B<3> ), .Cin(n17), .S(\S<3> ), .P(p3), .G(g3)
         );
  AND2X2 U1 ( .A(p1), .B(p0), .Y(n32) );
  AOI21X1 U12 ( .A(Cin), .B(P), .C(G), .Y(n35) );
  AOI21X1 U15 ( .A(g0), .B(p1), .C(g1), .Y(n34) );
  NAND3X1 U16 ( .A(p3), .B(p2), .C(n32), .Y(n33) );
  INVX1 U2 ( .A(g1), .Y(n24) );
  INVX1 U3 ( .A(g0), .Y(n23) );
  INVX1 U4 ( .A(g2), .Y(n22) );
  INVX1 U5 ( .A(p3), .Y(n28) );
  INVX1 U6 ( .A(g3), .Y(n27) );
  INVX1 U7 ( .A(n11), .Y(Cout) );
  AND2X1 U8 ( .A(Cin), .B(p0), .Y(n4) );
  AND2X2 U9 ( .A(p2), .B(n7), .Y(n2) );
  BUFX2 U10 ( .A(n20), .Y(n1) );
  INVX1 U11 ( .A(n2), .Y(n3) );
  INVX1 U13 ( .A(n4), .Y(n5) );
  AND2X2 U14 ( .A(n1), .B(n8), .Y(n6) );
  INVX1 U17 ( .A(n6), .Y(n7) );
  BUFX2 U18 ( .A(n21), .Y(n8) );
  BUFX2 U19 ( .A(n34), .Y(n9) );
  INVX1 U20 ( .A(n9), .Y(n26) );
  BUFX2 U21 ( .A(n35), .Y(n11) );
  INVX1 U22 ( .A(n33), .Y(P) );
  BUFX2 U23 ( .A(n29), .Y(n12) );
  AND2X2 U24 ( .A(n22), .B(n3), .Y(n16) );
  INVX1 U25 ( .A(n16), .Y(n17) );
  INVX1 U26 ( .A(n19), .Y(n18) );
  AND2X2 U27 ( .A(n5), .B(n23), .Y(n19) );
  AOI21X1 U28 ( .A(p1), .B(g0), .C(g1), .Y(n21) );
  NAND3X1 U29 ( .A(p1), .B(p0), .C(Cin), .Y(n20) );
  INVX2 U30 ( .A(p1), .Y(n25) );
  OAI21X1 U31 ( .A(n25), .B(n19), .C(n24), .Y(n30) );
  AOI21X1 U32 ( .A(n26), .B(p2), .C(g2), .Y(n29) );
  OAI21X1 U33 ( .A(n12), .B(n28), .C(n27), .Y(G) );
endmodule


module CLA4_7 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, Cout, P, G, .S({\S<3> , \S<2> , \S<1> , \S<0> }
        ) );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output Cout, P, G, \S<3> , \S<2> , \S<1> , \S<0> ;
  wire   p0, g0, p1, g1, p2, g2, c3, p3, g3, n1, n2, n3, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n23;

  pfa_31 bit0 ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(p0), .G(g0)
         );
  pfa_30 bit1 ( .A(\A<1> ), .B(\B<1> ), .Cin(n6), .S(\S<1> ), .P(p1), .G(g1)
         );
  pfa_29 bit2 ( .A(\A<2> ), .B(\B<2> ), .Cin(n23), .S(\S<2> ), .P(p2), .G(g2)
         );
  pfa_28 bit3 ( .A(\A<3> ), .B(\B<3> ), .Cin(c3), .S(\S<3> ), .P(p3), .G(g3)
         );
  INVX1 U1 ( .A(g2), .Y(n15) );
  INVX1 U2 ( .A(g1), .Y(n12) );
  INVX1 U3 ( .A(Cin), .Y(n20) );
  AND2X2 U4 ( .A(n18), .B(p3), .Y(n10) );
  OR2X2 U5 ( .A(g3), .B(n10), .Y(G) );
  AND2X2 U6 ( .A(Cin), .B(p0), .Y(n1) );
  INVX1 U7 ( .A(n1), .Y(n2) );
  BUFX2 U8 ( .A(n17), .Y(n3) );
  INVX1 U9 ( .A(G), .Y(n5) );
  INVX1 U10 ( .A(n7), .Y(n6) );
  AND2X2 U11 ( .A(n11), .B(n2), .Y(n7) );
  INVX1 U12 ( .A(P), .Y(n8) );
  BUFX2 U13 ( .A(n16), .Y(n9) );
  INVX1 U14 ( .A(n21), .Y(P) );
  INVX1 U15 ( .A(g0), .Y(n11) );
  INVX1 U16 ( .A(p2), .Y(n16) );
  INVX1 U17 ( .A(p1), .Y(n13) );
  OAI21X1 U18 ( .A(n7), .B(n13), .C(n12), .Y(n23) );
  INVX2 U19 ( .A(n23), .Y(n14) );
  OAI21X1 U20 ( .A(n9), .B(n14), .C(n15), .Y(c3) );
  AOI21X1 U21 ( .A(p1), .B(g0), .C(g1), .Y(n17) );
  OAI21X1 U22 ( .A(n16), .B(n3), .C(n15), .Y(n18) );
  AND2X2 U23 ( .A(p3), .B(p2), .Y(n19) );
  NAND3X1 U24 ( .A(p1), .B(p0), .C(n19), .Y(n21) );
  OAI21X1 U25 ( .A(n8), .B(n20), .C(n5), .Y(Cout) );
endmodule


module CLA4_6 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, Cout, P, G, .S({\S<3> , \S<2> , \S<1> , \S<0> }
        ) );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output Cout, P, G, \S<3> , \S<2> , \S<1> , \S<0> ;
  wire   p0, g0, p1, g1, p2, g2, p3, g3, n1, n2, n3, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n34;

  pfa_27 bit0 ( .A(\A<0> ), .B(\B<0> ), .Cin(n21), .S(\S<0> ), .P(p0), .G(g0)
         );
  pfa_26 bit1 ( .A(\A<1> ), .B(\B<1> ), .Cin(n2), .S(\S<1> ), .P(p1), .G(g1)
         );
  pfa_25 bit2 ( .A(\A<2> ), .B(\B<2> ), .Cin(n24), .S(\S<2> ), .P(p2), .G(g2)
         );
  pfa_24 bit3 ( .A(\A<3> ), .B(\B<3> ), .Cin(n14), .S(\S<3> ), .P(p3), .G(g3)
         );
  INVX1 U1 ( .A(g2), .Y(n27) );
  INVX1 U2 ( .A(p2), .Y(n28) );
  INVX1 U3 ( .A(g1), .Y(n25) );
  INVX1 U4 ( .A(g3), .Y(n31) );
  INVX1 U5 ( .A(p1), .Y(n26) );
  AND2X2 U6 ( .A(p2), .B(n34), .Y(n10) );
  AND2X2 U7 ( .A(n21), .B(P), .Y(n11) );
  AND2X2 U8 ( .A(n22), .B(n20), .Y(n1) );
  INVX1 U9 ( .A(n1), .Y(n2) );
  AND2X2 U10 ( .A(n31), .B(n6), .Y(n3) );
  INVX1 U11 ( .A(n3), .Y(G) );
  AND2X2 U12 ( .A(p3), .B(n30), .Y(n5) );
  INVX1 U13 ( .A(n5), .Y(n6) );
  BUFX2 U14 ( .A(n32), .Y(n7) );
  BUFX2 U15 ( .A(n29), .Y(n8) );
  INVX1 U16 ( .A(n10), .Y(n9) );
  INVX1 U17 ( .A(n11), .Y(n12) );
  AND2X2 U18 ( .A(n27), .B(n9), .Y(n13) );
  INVX1 U19 ( .A(n13), .Y(n14) );
  AND2X2 U20 ( .A(Cin), .B(p0), .Y(n15) );
  INVX1 U21 ( .A(n15), .Y(n16) );
  OR2X2 U22 ( .A(n7), .B(n26), .Y(n17) );
  INVX1 U23 ( .A(n17), .Y(P) );
  INVX1 U24 ( .A(n16), .Y(n19) );
  INVX1 U25 ( .A(n19), .Y(n20) );
  INVX1 U26 ( .A(g0), .Y(n22) );
  BUFX2 U27 ( .A(Cin), .Y(n21) );
  AND2X2 U28 ( .A(n16), .B(n22), .Y(n23) );
  OAI21X1 U29 ( .A(n23), .B(n26), .C(n25), .Y(n24) );
  OAI21X1 U30 ( .A(n23), .B(n26), .C(n25), .Y(n34) );
  AOI21X1 U31 ( .A(p1), .B(g0), .C(g1), .Y(n29) );
  OAI21X1 U32 ( .A(n8), .B(n28), .C(n27), .Y(n30) );
  NAND3X1 U33 ( .A(p3), .B(p2), .C(p0), .Y(n32) );
  NAND2X1 U34 ( .A(n3), .B(n12), .Y(Cout) );
endmodule


module CLA4_5 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, Cout, P, G, .S({\S<3> , \S<2> , \S<1> , \S<0> }
        ) );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output Cout, P, G, \S<3> , \S<2> , \S<1> , \S<0> ;
  wire   p0, g0, p1, g1, p2, g2, p3, g3, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n21, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n33;

  pfa_23 bit0 ( .A(\A<0> ), .B(\B<0> ), .Cin(n1), .S(\S<0> ), .P(p0), .G(g0)
         );
  pfa_22 bit1 ( .A(\A<1> ), .B(\B<1> ), .Cin(n4), .S(\S<1> ), .P(p1), .G(g1)
         );
  pfa_21 bit2 ( .A(\A<2> ), .B(\B<2> ), .Cin(n3), .S(\S<2> ), .P(p2), .G(g2)
         );
  pfa_20 bit3 ( .A(\A<3> ), .B(\B<3> ), .Cin(n18), .S(\S<3> ), .P(p3), .G(g3)
         );
  INVX1 U1 ( .A(p2), .Y(n26) );
  INVX1 U2 ( .A(g0), .Y(n24) );
  INVX1 U3 ( .A(g2), .Y(n25) );
  INVX1 U4 ( .A(p1), .Y(n31) );
  INVX1 U5 ( .A(g3), .Y(n29) );
  BUFX2 U6 ( .A(Cin), .Y(n1) );
  INVX1 U7 ( .A(n33), .Y(n2) );
  INVX1 U8 ( .A(n2), .Y(n3) );
  AND2X1 U9 ( .A(Cin), .B(p0), .Y(n5) );
  AND2X2 U10 ( .A(p2), .B(n33), .Y(n8) );
  INVX1 U11 ( .A(n7), .Y(n4) );
  AND2X2 U12 ( .A(n24), .B(n6), .Y(n7) );
  INVX1 U13 ( .A(n5), .Y(n6) );
  INVX1 U14 ( .A(n8), .Y(n9) );
  AND2X2 U15 ( .A(p3), .B(n28), .Y(n10) );
  INVX1 U16 ( .A(n10), .Y(n11) );
  AND2X1 U17 ( .A(n1), .B(P), .Y(n12) );
  INVX1 U18 ( .A(n12), .Y(n13) );
  INVX1 U19 ( .A(n30), .Y(n14) );
  INVX1 U20 ( .A(n14), .Y(n15) );
  INVX1 U21 ( .A(n23), .Y(n33) );
  BUFX2 U22 ( .A(n27), .Y(n16) );
  AND2X2 U23 ( .A(n25), .B(n9), .Y(n17) );
  INVX1 U24 ( .A(n17), .Y(n18) );
  OR2X2 U25 ( .A(n31), .B(n15), .Y(n19) );
  INVX1 U26 ( .A(n19), .Y(P) );
  AND2X2 U27 ( .A(n29), .B(n11), .Y(n21) );
  INVX1 U28 ( .A(n21), .Y(G) );
  AOI21X1 U29 ( .A(n4), .B(p1), .C(g1), .Y(n23) );
  AOI21X1 U30 ( .A(p1), .B(g0), .C(g1), .Y(n27) );
  OAI21X1 U31 ( .A(n16), .B(n26), .C(n25), .Y(n28) );
  NAND3X1 U32 ( .A(p3), .B(p2), .C(p0), .Y(n30) );
  NAND2X1 U33 ( .A(n21), .B(n13), .Y(Cout) );
endmodule


module CLA4_4 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, Cout, P, G, .S({\S<3> , \S<2> , \S<1> , \S<0> }
        ) );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output Cout, P, G, \S<3> , \S<2> , \S<1> , \S<0> ;
  wire   p0, g0, p1, g1, p2, g2, p3, g3, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32;

  pfa_19 bit0 ( .A(\A<0> ), .B(\B<0> ), .Cin(n23), .S(\S<0> ), .P(p0), .G(g0)
         );
  pfa_18 bit1 ( .A(\A<1> ), .B(\B<1> ), .Cin(n19), .S(\S<1> ), .P(p1), .G(g1)
         );
  pfa_17 bit2 ( .A(\A<2> ), .B(\B<2> ), .Cin(n18), .S(\S<2> ), .P(p2), .G(g2)
         );
  pfa_16 bit3 ( .A(\A<3> ), .B(\B<3> ), .Cin(n16), .S(\S<3> ), .P(p3), .G(g3)
         );
  AOI21X1 U12 ( .A(n23), .B(P), .C(G), .Y(n32) );
  AOI21X1 U13 ( .A(p3), .B(n30), .C(g3), .Y(n31) );
  OAI21X1 U14 ( .A(n9), .B(n25), .C(n26), .Y(n30) );
  AOI21X1 U15 ( .A(g0), .B(p1), .C(g1), .Y(n29) );
  NAND3X1 U16 ( .A(p3), .B(p2), .C(n27), .Y(n28) );
  INVX1 U1 ( .A(g1), .Y(n24) );
  INVX1 U2 ( .A(p2), .Y(n25) );
  INVX1 U3 ( .A(g2), .Y(n26) );
  BUFX2 U4 ( .A(Cin), .Y(n23) );
  OR2X2 U5 ( .A(n3), .B(g0), .Y(n1) );
  INVX1 U6 ( .A(n1), .Y(n20) );
  INVX2 U7 ( .A(n2), .Y(n16) );
  OAI21X1 U8 ( .A(n8), .B(n22), .C(n4), .Y(n2) );
  AND2X2 U9 ( .A(n24), .B(n21), .Y(n17) );
  AND2X2 U10 ( .A(p0), .B(Cin), .Y(n3) );
  AND2X1 U11 ( .A(p1), .B(p0), .Y(n27) );
  OR2X1 U17 ( .A(g2), .B(p2), .Y(n4) );
  BUFX2 U18 ( .A(n28), .Y(n5) );
  INVX1 U19 ( .A(n5), .Y(P) );
  BUFX2 U20 ( .A(n31), .Y(n6) );
  INVX1 U21 ( .A(n6), .Y(G) );
  BUFX2 U22 ( .A(n32), .Y(n7) );
  INVX1 U23 ( .A(n7), .Y(Cout) );
  OR2X1 U24 ( .A(g1), .B(g2), .Y(n8) );
  BUFX2 U25 ( .A(n29), .Y(n9) );
  INVX1 U26 ( .A(n17), .Y(n18) );
  INVX1 U27 ( .A(n20), .Y(n19) );
  INVX1 U28 ( .A(n22), .Y(n21) );
  AND2X2 U29 ( .A(n1), .B(p1), .Y(n22) );
endmodule


module reg16_7 ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n1, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84;

  dff_127 d0 ( .q(\read<0> ), .d(n84), .clk(clk), .rst(rst) );
  dff_126 d1 ( .q(\read<1> ), .d(n83), .clk(clk), .rst(rst) );
  dff_125 d2 ( .q(\read<2> ), .d(n82), .clk(clk), .rst(rst) );
  dff_124 d3 ( .q(\read<3> ), .d(n81), .clk(clk), .rst(rst) );
  dff_123 d4 ( .q(\read<4> ), .d(n80), .clk(clk), .rst(rst) );
  dff_122 d5 ( .q(\read<5> ), .d(n79), .clk(clk), .rst(rst) );
  dff_121 d6 ( .q(\read<6> ), .d(n78), .clk(clk), .rst(rst) );
  dff_120 d7 ( .q(\read<7> ), .d(n77), .clk(clk), .rst(rst) );
  dff_119 d8 ( .q(\read<8> ), .d(n76), .clk(clk), .rst(rst) );
  dff_118 d9 ( .q(\read<9> ), .d(n75), .clk(clk), .rst(rst) );
  dff_117 d10 ( .q(\read<10> ), .d(n74), .clk(clk), .rst(rst) );
  dff_116 d11 ( .q(\read<11> ), .d(n73), .clk(clk), .rst(rst) );
  dff_115 d12 ( .q(\read<12> ), .d(n72), .clk(clk), .rst(rst) );
  dff_114 d13 ( .q(\read<13> ), .d(n71), .clk(clk), .rst(rst) );
  dff_113 d14 ( .q(\read<14> ), .d(n70), .clk(clk), .rst(rst) );
  dff_112 d15 ( .q(\read<15> ), .d(n69), .clk(clk), .rst(rst) );
  AOI22X1 U18 ( .A(\read<9> ), .B(n68), .C(\write<9> ), .D(n50), .Y(n67) );
  AOI22X1 U19 ( .A(\read<8> ), .B(n68), .C(\write<8> ), .D(n50), .Y(n66) );
  AOI22X1 U20 ( .A(\read<7> ), .B(n68), .C(\write<7> ), .D(n50), .Y(n65) );
  AOI22X1 U21 ( .A(\read<6> ), .B(n68), .C(\write<6> ), .D(n50), .Y(n64) );
  AOI22X1 U22 ( .A(\read<5> ), .B(n68), .C(\write<5> ), .D(n50), .Y(n63) );
  AOI22X1 U23 ( .A(\read<4> ), .B(n68), .C(\write<4> ), .D(n50), .Y(n62) );
  AOI22X1 U24 ( .A(\read<3> ), .B(n68), .C(\write<3> ), .D(n51), .Y(n61) );
  AOI22X1 U25 ( .A(\read<2> ), .B(n68), .C(\write<2> ), .D(n51), .Y(n60) );
  AOI22X1 U26 ( .A(\read<1> ), .B(n68), .C(\write<1> ), .D(n51), .Y(n59) );
  AOI22X1 U27 ( .A(\read<15> ), .B(n68), .C(\write<15> ), .D(n51), .Y(n58) );
  AOI22X1 U28 ( .A(\read<14> ), .B(n68), .C(\write<14> ), .D(n51), .Y(n57) );
  AOI22X1 U29 ( .A(\read<13> ), .B(n68), .C(\write<13> ), .D(n51), .Y(n56) );
  AOI22X1 U30 ( .A(\read<12> ), .B(n68), .C(\write<12> ), .D(n51), .Y(n55) );
  AOI22X1 U31 ( .A(\read<11> ), .B(n68), .C(\write<11> ), .D(n51), .Y(n54) );
  AOI22X1 U32 ( .A(\read<10> ), .B(n68), .C(\write<10> ), .D(n51), .Y(n53) );
  AOI22X1 U33 ( .A(\read<0> ), .B(n68), .C(\write<0> ), .D(n51), .Y(n52) );
  BUFX2 U1 ( .A(wr_en), .Y(n50) );
  BUFX2 U2 ( .A(wr_en), .Y(n51) );
  INVX1 U3 ( .A(n50), .Y(n68) );
  BUFX2 U4 ( .A(n52), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n84) );
  BUFX2 U6 ( .A(n53), .Y(n35) );
  INVX1 U7 ( .A(n35), .Y(n74) );
  BUFX2 U8 ( .A(n54), .Y(n36) );
  INVX1 U9 ( .A(n36), .Y(n73) );
  BUFX2 U10 ( .A(n55), .Y(n37) );
  INVX1 U11 ( .A(n37), .Y(n72) );
  BUFX2 U12 ( .A(n56), .Y(n38) );
  INVX1 U13 ( .A(n38), .Y(n71) );
  BUFX2 U14 ( .A(n57), .Y(n39) );
  INVX1 U15 ( .A(n39), .Y(n70) );
  BUFX2 U16 ( .A(n58), .Y(n40) );
  INVX1 U17 ( .A(n40), .Y(n69) );
  BUFX2 U34 ( .A(n59), .Y(n41) );
  INVX1 U35 ( .A(n41), .Y(n83) );
  BUFX2 U36 ( .A(n60), .Y(n42) );
  INVX1 U37 ( .A(n42), .Y(n82) );
  BUFX2 U38 ( .A(n61), .Y(n43) );
  INVX1 U39 ( .A(n43), .Y(n81) );
  BUFX2 U40 ( .A(n62), .Y(n44) );
  INVX1 U41 ( .A(n44), .Y(n80) );
  BUFX2 U42 ( .A(n63), .Y(n45) );
  INVX1 U43 ( .A(n45), .Y(n79) );
  BUFX2 U44 ( .A(n64), .Y(n46) );
  INVX1 U45 ( .A(n46), .Y(n78) );
  BUFX2 U46 ( .A(n65), .Y(n47) );
  INVX1 U47 ( .A(n47), .Y(n77) );
  BUFX2 U48 ( .A(n66), .Y(n48) );
  INVX1 U49 ( .A(n48), .Y(n76) );
  BUFX2 U50 ( .A(n67), .Y(n49) );
  INVX1 U51 ( .A(n49), .Y(n75) );
endmodule


module reg16_6 ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n1, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84;

  dff_111 d0 ( .q(\read<0> ), .d(n84), .clk(clk), .rst(rst) );
  dff_110 d1 ( .q(\read<1> ), .d(n83), .clk(clk), .rst(rst) );
  dff_109 d2 ( .q(\read<2> ), .d(n82), .clk(clk), .rst(rst) );
  dff_108 d3 ( .q(\read<3> ), .d(n81), .clk(clk), .rst(rst) );
  dff_107 d4 ( .q(\read<4> ), .d(n80), .clk(clk), .rst(rst) );
  dff_106 d5 ( .q(\read<5> ), .d(n79), .clk(clk), .rst(rst) );
  dff_105 d6 ( .q(\read<6> ), .d(n78), .clk(clk), .rst(rst) );
  dff_104 d7 ( .q(\read<7> ), .d(n77), .clk(clk), .rst(rst) );
  dff_103 d8 ( .q(\read<8> ), .d(n76), .clk(clk), .rst(rst) );
  dff_102 d9 ( .q(\read<9> ), .d(n75), .clk(clk), .rst(rst) );
  dff_101 d10 ( .q(\read<10> ), .d(n74), .clk(clk), .rst(rst) );
  dff_100 d11 ( .q(\read<11> ), .d(n73), .clk(clk), .rst(rst) );
  dff_99 d12 ( .q(\read<12> ), .d(n72), .clk(clk), .rst(rst) );
  dff_98 d13 ( .q(\read<13> ), .d(n71), .clk(clk), .rst(rst) );
  dff_97 d14 ( .q(\read<14> ), .d(n70), .clk(clk), .rst(rst) );
  dff_96 d15 ( .q(\read<15> ), .d(n69), .clk(clk), .rst(rst) );
  AOI22X1 U18 ( .A(\read<9> ), .B(n68), .C(\write<9> ), .D(n50), .Y(n67) );
  AOI22X1 U19 ( .A(\read<8> ), .B(n68), .C(\write<8> ), .D(n50), .Y(n66) );
  AOI22X1 U20 ( .A(\read<7> ), .B(n68), .C(\write<7> ), .D(n50), .Y(n65) );
  AOI22X1 U21 ( .A(\read<6> ), .B(n68), .C(\write<6> ), .D(n50), .Y(n64) );
  AOI22X1 U22 ( .A(\read<5> ), .B(n68), .C(\write<5> ), .D(n50), .Y(n63) );
  AOI22X1 U23 ( .A(\read<4> ), .B(n68), .C(\write<4> ), .D(n50), .Y(n62) );
  AOI22X1 U24 ( .A(\read<3> ), .B(n68), .C(\write<3> ), .D(n51), .Y(n61) );
  AOI22X1 U25 ( .A(\read<2> ), .B(n68), .C(\write<2> ), .D(n51), .Y(n60) );
  AOI22X1 U26 ( .A(\read<1> ), .B(n68), .C(\write<1> ), .D(n51), .Y(n59) );
  AOI22X1 U27 ( .A(\read<15> ), .B(n68), .C(\write<15> ), .D(n51), .Y(n58) );
  AOI22X1 U28 ( .A(\read<14> ), .B(n68), .C(\write<14> ), .D(n51), .Y(n57) );
  AOI22X1 U29 ( .A(\read<13> ), .B(n68), .C(\write<13> ), .D(n51), .Y(n56) );
  AOI22X1 U30 ( .A(\read<12> ), .B(n68), .C(\write<12> ), .D(n51), .Y(n55) );
  AOI22X1 U31 ( .A(\read<11> ), .B(n68), .C(\write<11> ), .D(n51), .Y(n54) );
  AOI22X1 U32 ( .A(\read<10> ), .B(n68), .C(\write<10> ), .D(n51), .Y(n53) );
  AOI22X1 U33 ( .A(\read<0> ), .B(n68), .C(\write<0> ), .D(n51), .Y(n52) );
  BUFX2 U1 ( .A(wr_en), .Y(n50) );
  BUFX2 U2 ( .A(wr_en), .Y(n51) );
  INVX1 U3 ( .A(n50), .Y(n68) );
  BUFX2 U4 ( .A(n52), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n84) );
  BUFX2 U6 ( .A(n53), .Y(n35) );
  INVX1 U7 ( .A(n35), .Y(n74) );
  BUFX2 U8 ( .A(n54), .Y(n36) );
  INVX1 U9 ( .A(n36), .Y(n73) );
  BUFX2 U10 ( .A(n55), .Y(n37) );
  INVX1 U11 ( .A(n37), .Y(n72) );
  BUFX2 U12 ( .A(n56), .Y(n38) );
  INVX1 U13 ( .A(n38), .Y(n71) );
  BUFX2 U14 ( .A(n57), .Y(n39) );
  INVX1 U15 ( .A(n39), .Y(n70) );
  BUFX2 U16 ( .A(n58), .Y(n40) );
  INVX1 U17 ( .A(n40), .Y(n69) );
  BUFX2 U34 ( .A(n59), .Y(n41) );
  INVX1 U35 ( .A(n41), .Y(n83) );
  BUFX2 U36 ( .A(n60), .Y(n42) );
  INVX1 U37 ( .A(n42), .Y(n82) );
  BUFX2 U38 ( .A(n61), .Y(n43) );
  INVX1 U39 ( .A(n43), .Y(n81) );
  BUFX2 U40 ( .A(n62), .Y(n44) );
  INVX1 U41 ( .A(n44), .Y(n80) );
  BUFX2 U42 ( .A(n63), .Y(n45) );
  INVX1 U43 ( .A(n45), .Y(n79) );
  BUFX2 U44 ( .A(n64), .Y(n46) );
  INVX1 U45 ( .A(n46), .Y(n78) );
  BUFX2 U46 ( .A(n65), .Y(n47) );
  INVX1 U47 ( .A(n47), .Y(n77) );
  BUFX2 U48 ( .A(n66), .Y(n48) );
  INVX1 U49 ( .A(n48), .Y(n76) );
  BUFX2 U50 ( .A(n67), .Y(n49) );
  INVX1 U51 ( .A(n49), .Y(n75) );
endmodule


module reg16_5 ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n1, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84;

  dff_95 d0 ( .q(\read<0> ), .d(n84), .clk(clk), .rst(rst) );
  dff_94 d1 ( .q(\read<1> ), .d(n83), .clk(clk), .rst(rst) );
  dff_93 d2 ( .q(\read<2> ), .d(n82), .clk(clk), .rst(rst) );
  dff_92 d3 ( .q(\read<3> ), .d(n81), .clk(clk), .rst(rst) );
  dff_91 d4 ( .q(\read<4> ), .d(n80), .clk(clk), .rst(rst) );
  dff_90 d5 ( .q(\read<5> ), .d(n79), .clk(clk), .rst(rst) );
  dff_89 d6 ( .q(\read<6> ), .d(n78), .clk(clk), .rst(rst) );
  dff_88 d7 ( .q(\read<7> ), .d(n77), .clk(clk), .rst(rst) );
  dff_87 d8 ( .q(\read<8> ), .d(n76), .clk(clk), .rst(rst) );
  dff_86 d9 ( .q(\read<9> ), .d(n75), .clk(clk), .rst(rst) );
  dff_85 d10 ( .q(\read<10> ), .d(n74), .clk(clk), .rst(rst) );
  dff_84 d11 ( .q(\read<11> ), .d(n73), .clk(clk), .rst(rst) );
  dff_83 d12 ( .q(\read<12> ), .d(n72), .clk(clk), .rst(rst) );
  dff_82 d13 ( .q(\read<13> ), .d(n71), .clk(clk), .rst(rst) );
  dff_81 d14 ( .q(\read<14> ), .d(n70), .clk(clk), .rst(rst) );
  dff_80 d15 ( .q(\read<15> ), .d(n69), .clk(clk), .rst(rst) );
  AOI22X1 U18 ( .A(\read<9> ), .B(n68), .C(\write<9> ), .D(n50), .Y(n67) );
  AOI22X1 U19 ( .A(\read<8> ), .B(n68), .C(\write<8> ), .D(n50), .Y(n66) );
  AOI22X1 U20 ( .A(\read<7> ), .B(n68), .C(\write<7> ), .D(n50), .Y(n65) );
  AOI22X1 U21 ( .A(\read<6> ), .B(n68), .C(\write<6> ), .D(n50), .Y(n64) );
  AOI22X1 U22 ( .A(\read<5> ), .B(n68), .C(\write<5> ), .D(n50), .Y(n63) );
  AOI22X1 U23 ( .A(\read<4> ), .B(n68), .C(\write<4> ), .D(n50), .Y(n62) );
  AOI22X1 U24 ( .A(\read<3> ), .B(n68), .C(\write<3> ), .D(n51), .Y(n61) );
  AOI22X1 U25 ( .A(\read<2> ), .B(n68), .C(\write<2> ), .D(n51), .Y(n60) );
  AOI22X1 U26 ( .A(\read<1> ), .B(n68), .C(\write<1> ), .D(n51), .Y(n59) );
  AOI22X1 U27 ( .A(\read<15> ), .B(n68), .C(\write<15> ), .D(n51), .Y(n58) );
  AOI22X1 U28 ( .A(\read<14> ), .B(n68), .C(\write<14> ), .D(n51), .Y(n57) );
  AOI22X1 U29 ( .A(\read<13> ), .B(n68), .C(\write<13> ), .D(n51), .Y(n56) );
  AOI22X1 U30 ( .A(\read<12> ), .B(n68), .C(\write<12> ), .D(n51), .Y(n55) );
  AOI22X1 U31 ( .A(\read<11> ), .B(n68), .C(\write<11> ), .D(n51), .Y(n54) );
  AOI22X1 U32 ( .A(\read<10> ), .B(n68), .C(\write<10> ), .D(n51), .Y(n53) );
  AOI22X1 U33 ( .A(\read<0> ), .B(n68), .C(\write<0> ), .D(n51), .Y(n52) );
  BUFX2 U1 ( .A(wr_en), .Y(n50) );
  BUFX2 U2 ( .A(wr_en), .Y(n51) );
  INVX1 U3 ( .A(n50), .Y(n68) );
  BUFX2 U4 ( .A(n52), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n84) );
  BUFX2 U6 ( .A(n53), .Y(n35) );
  INVX1 U7 ( .A(n35), .Y(n74) );
  BUFX2 U8 ( .A(n54), .Y(n36) );
  INVX1 U9 ( .A(n36), .Y(n73) );
  BUFX2 U10 ( .A(n55), .Y(n37) );
  INVX1 U11 ( .A(n37), .Y(n72) );
  BUFX2 U12 ( .A(n56), .Y(n38) );
  INVX1 U13 ( .A(n38), .Y(n71) );
  BUFX2 U14 ( .A(n57), .Y(n39) );
  INVX1 U15 ( .A(n39), .Y(n70) );
  BUFX2 U16 ( .A(n58), .Y(n40) );
  INVX1 U17 ( .A(n40), .Y(n69) );
  BUFX2 U34 ( .A(n59), .Y(n41) );
  INVX1 U35 ( .A(n41), .Y(n83) );
  BUFX2 U36 ( .A(n60), .Y(n42) );
  INVX1 U37 ( .A(n42), .Y(n82) );
  BUFX2 U38 ( .A(n61), .Y(n43) );
  INVX1 U39 ( .A(n43), .Y(n81) );
  BUFX2 U40 ( .A(n62), .Y(n44) );
  INVX1 U41 ( .A(n44), .Y(n80) );
  BUFX2 U42 ( .A(n63), .Y(n45) );
  INVX1 U43 ( .A(n45), .Y(n79) );
  BUFX2 U44 ( .A(n64), .Y(n46) );
  INVX1 U45 ( .A(n46), .Y(n78) );
  BUFX2 U46 ( .A(n65), .Y(n47) );
  INVX1 U47 ( .A(n47), .Y(n77) );
  BUFX2 U48 ( .A(n66), .Y(n48) );
  INVX1 U49 ( .A(n48), .Y(n76) );
  BUFX2 U50 ( .A(n67), .Y(n49) );
  INVX1 U51 ( .A(n49), .Y(n75) );
endmodule


module reg16_4 ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n1, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84;

  dff_79 d0 ( .q(\read<0> ), .d(n84), .clk(clk), .rst(rst) );
  dff_78 d1 ( .q(\read<1> ), .d(n83), .clk(clk), .rst(rst) );
  dff_77 d2 ( .q(\read<2> ), .d(n82), .clk(clk), .rst(rst) );
  dff_76 d3 ( .q(\read<3> ), .d(n81), .clk(clk), .rst(rst) );
  dff_75 d4 ( .q(\read<4> ), .d(n80), .clk(clk), .rst(rst) );
  dff_74 d5 ( .q(\read<5> ), .d(n79), .clk(clk), .rst(rst) );
  dff_73 d6 ( .q(\read<6> ), .d(n78), .clk(clk), .rst(rst) );
  dff_72 d7 ( .q(\read<7> ), .d(n77), .clk(clk), .rst(rst) );
  dff_71 d8 ( .q(\read<8> ), .d(n76), .clk(clk), .rst(rst) );
  dff_70 d9 ( .q(\read<9> ), .d(n75), .clk(clk), .rst(rst) );
  dff_69 d10 ( .q(\read<10> ), .d(n74), .clk(clk), .rst(rst) );
  dff_68 d11 ( .q(\read<11> ), .d(n73), .clk(clk), .rst(rst) );
  dff_67 d12 ( .q(\read<12> ), .d(n72), .clk(clk), .rst(rst) );
  dff_66 d13 ( .q(\read<13> ), .d(n71), .clk(clk), .rst(rst) );
  dff_65 d14 ( .q(\read<14> ), .d(n70), .clk(clk), .rst(rst) );
  dff_64 d15 ( .q(\read<15> ), .d(n69), .clk(clk), .rst(rst) );
  AOI22X1 U18 ( .A(\read<9> ), .B(n68), .C(\write<9> ), .D(n50), .Y(n67) );
  AOI22X1 U19 ( .A(\read<8> ), .B(n68), .C(\write<8> ), .D(n50), .Y(n66) );
  AOI22X1 U20 ( .A(\read<7> ), .B(n68), .C(\write<7> ), .D(n50), .Y(n65) );
  AOI22X1 U21 ( .A(\read<6> ), .B(n68), .C(\write<6> ), .D(n50), .Y(n64) );
  AOI22X1 U22 ( .A(\read<5> ), .B(n68), .C(\write<5> ), .D(n50), .Y(n63) );
  AOI22X1 U23 ( .A(\read<4> ), .B(n68), .C(\write<4> ), .D(n50), .Y(n62) );
  AOI22X1 U24 ( .A(\read<3> ), .B(n68), .C(\write<3> ), .D(n51), .Y(n61) );
  AOI22X1 U25 ( .A(\read<2> ), .B(n68), .C(\write<2> ), .D(n51), .Y(n60) );
  AOI22X1 U26 ( .A(\read<1> ), .B(n68), .C(\write<1> ), .D(n51), .Y(n59) );
  AOI22X1 U27 ( .A(\read<15> ), .B(n68), .C(\write<15> ), .D(n51), .Y(n58) );
  AOI22X1 U28 ( .A(\read<14> ), .B(n68), .C(\write<14> ), .D(n51), .Y(n57) );
  AOI22X1 U29 ( .A(\read<13> ), .B(n68), .C(\write<13> ), .D(n51), .Y(n56) );
  AOI22X1 U30 ( .A(\read<12> ), .B(n68), .C(\write<12> ), .D(n51), .Y(n55) );
  AOI22X1 U31 ( .A(\read<11> ), .B(n68), .C(\write<11> ), .D(n51), .Y(n54) );
  AOI22X1 U32 ( .A(\read<10> ), .B(n68), .C(\write<10> ), .D(n51), .Y(n53) );
  AOI22X1 U33 ( .A(\read<0> ), .B(n68), .C(\write<0> ), .D(n51), .Y(n52) );
  BUFX2 U1 ( .A(wr_en), .Y(n50) );
  BUFX2 U2 ( .A(wr_en), .Y(n51) );
  INVX1 U3 ( .A(n50), .Y(n68) );
  BUFX2 U4 ( .A(n52), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n84) );
  BUFX2 U6 ( .A(n53), .Y(n35) );
  INVX1 U7 ( .A(n35), .Y(n74) );
  BUFX2 U8 ( .A(n54), .Y(n36) );
  INVX1 U9 ( .A(n36), .Y(n73) );
  BUFX2 U10 ( .A(n55), .Y(n37) );
  INVX1 U11 ( .A(n37), .Y(n72) );
  BUFX2 U12 ( .A(n56), .Y(n38) );
  INVX1 U13 ( .A(n38), .Y(n71) );
  BUFX2 U14 ( .A(n57), .Y(n39) );
  INVX1 U15 ( .A(n39), .Y(n70) );
  BUFX2 U16 ( .A(n58), .Y(n40) );
  INVX1 U17 ( .A(n40), .Y(n69) );
  BUFX2 U34 ( .A(n59), .Y(n41) );
  INVX1 U35 ( .A(n41), .Y(n83) );
  BUFX2 U36 ( .A(n60), .Y(n42) );
  INVX1 U37 ( .A(n42), .Y(n82) );
  BUFX2 U38 ( .A(n61), .Y(n43) );
  INVX1 U39 ( .A(n43), .Y(n81) );
  BUFX2 U40 ( .A(n62), .Y(n44) );
  INVX1 U41 ( .A(n44), .Y(n80) );
  BUFX2 U42 ( .A(n63), .Y(n45) );
  INVX1 U43 ( .A(n45), .Y(n79) );
  BUFX2 U44 ( .A(n64), .Y(n46) );
  INVX1 U45 ( .A(n46), .Y(n78) );
  BUFX2 U46 ( .A(n65), .Y(n47) );
  INVX1 U47 ( .A(n47), .Y(n77) );
  BUFX2 U48 ( .A(n66), .Y(n48) );
  INVX1 U49 ( .A(n48), .Y(n76) );
  BUFX2 U50 ( .A(n67), .Y(n49) );
  INVX1 U51 ( .A(n49), .Y(n75) );
endmodule


module reg16_3 ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n1, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84;

  dff_63 d0 ( .q(\read<0> ), .d(n84), .clk(clk), .rst(rst) );
  dff_62 d1 ( .q(\read<1> ), .d(n83), .clk(clk), .rst(rst) );
  dff_61 d2 ( .q(\read<2> ), .d(n82), .clk(clk), .rst(rst) );
  dff_60 d3 ( .q(\read<3> ), .d(n81), .clk(clk), .rst(rst) );
  dff_59 d4 ( .q(\read<4> ), .d(n80), .clk(clk), .rst(rst) );
  dff_58 d5 ( .q(\read<5> ), .d(n79), .clk(clk), .rst(rst) );
  dff_57 d6 ( .q(\read<6> ), .d(n78), .clk(clk), .rst(rst) );
  dff_56 d7 ( .q(\read<7> ), .d(n77), .clk(clk), .rst(rst) );
  dff_55 d8 ( .q(\read<8> ), .d(n76), .clk(clk), .rst(rst) );
  dff_54 d9 ( .q(\read<9> ), .d(n75), .clk(clk), .rst(rst) );
  dff_53 d10 ( .q(\read<10> ), .d(n74), .clk(clk), .rst(rst) );
  dff_52 d11 ( .q(\read<11> ), .d(n73), .clk(clk), .rst(rst) );
  dff_51 d12 ( .q(\read<12> ), .d(n72), .clk(clk), .rst(rst) );
  dff_50 d13 ( .q(\read<13> ), .d(n71), .clk(clk), .rst(rst) );
  dff_49 d14 ( .q(\read<14> ), .d(n70), .clk(clk), .rst(rst) );
  dff_48 d15 ( .q(\read<15> ), .d(n69), .clk(clk), .rst(rst) );
  AOI22X1 U18 ( .A(\read<9> ), .B(n68), .C(\write<9> ), .D(n50), .Y(n67) );
  AOI22X1 U19 ( .A(\read<8> ), .B(n68), .C(\write<8> ), .D(n50), .Y(n66) );
  AOI22X1 U20 ( .A(\read<7> ), .B(n68), .C(\write<7> ), .D(n50), .Y(n65) );
  AOI22X1 U21 ( .A(\read<6> ), .B(n68), .C(\write<6> ), .D(n50), .Y(n64) );
  AOI22X1 U22 ( .A(\read<5> ), .B(n68), .C(\write<5> ), .D(n50), .Y(n63) );
  AOI22X1 U23 ( .A(\read<4> ), .B(n68), .C(\write<4> ), .D(n50), .Y(n62) );
  AOI22X1 U24 ( .A(\read<3> ), .B(n68), .C(\write<3> ), .D(n51), .Y(n61) );
  AOI22X1 U25 ( .A(\read<2> ), .B(n68), .C(\write<2> ), .D(n51), .Y(n60) );
  AOI22X1 U26 ( .A(\read<1> ), .B(n68), .C(\write<1> ), .D(n51), .Y(n59) );
  AOI22X1 U27 ( .A(\read<15> ), .B(n68), .C(\write<15> ), .D(n51), .Y(n58) );
  AOI22X1 U28 ( .A(\read<14> ), .B(n68), .C(\write<14> ), .D(n51), .Y(n57) );
  AOI22X1 U29 ( .A(\read<13> ), .B(n68), .C(\write<13> ), .D(n51), .Y(n56) );
  AOI22X1 U30 ( .A(\read<12> ), .B(n68), .C(\write<12> ), .D(n51), .Y(n55) );
  AOI22X1 U31 ( .A(\read<11> ), .B(n68), .C(\write<11> ), .D(n51), .Y(n54) );
  AOI22X1 U32 ( .A(\read<10> ), .B(n68), .C(\write<10> ), .D(n51), .Y(n53) );
  AOI22X1 U33 ( .A(\read<0> ), .B(n68), .C(\write<0> ), .D(n51), .Y(n52) );
  BUFX2 U1 ( .A(wr_en), .Y(n50) );
  BUFX2 U2 ( .A(wr_en), .Y(n51) );
  INVX1 U3 ( .A(n50), .Y(n68) );
  BUFX2 U4 ( .A(n52), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n84) );
  BUFX2 U6 ( .A(n53), .Y(n35) );
  INVX1 U7 ( .A(n35), .Y(n74) );
  BUFX2 U8 ( .A(n54), .Y(n36) );
  INVX1 U9 ( .A(n36), .Y(n73) );
  BUFX2 U10 ( .A(n55), .Y(n37) );
  INVX1 U11 ( .A(n37), .Y(n72) );
  BUFX2 U12 ( .A(n56), .Y(n38) );
  INVX1 U13 ( .A(n38), .Y(n71) );
  BUFX2 U14 ( .A(n57), .Y(n39) );
  INVX1 U15 ( .A(n39), .Y(n70) );
  BUFX2 U16 ( .A(n58), .Y(n40) );
  INVX1 U17 ( .A(n40), .Y(n69) );
  BUFX2 U34 ( .A(n59), .Y(n41) );
  INVX1 U35 ( .A(n41), .Y(n83) );
  BUFX2 U36 ( .A(n60), .Y(n42) );
  INVX1 U37 ( .A(n42), .Y(n82) );
  BUFX2 U38 ( .A(n61), .Y(n43) );
  INVX1 U39 ( .A(n43), .Y(n81) );
  BUFX2 U40 ( .A(n62), .Y(n44) );
  INVX1 U41 ( .A(n44), .Y(n80) );
  BUFX2 U42 ( .A(n63), .Y(n45) );
  INVX1 U43 ( .A(n45), .Y(n79) );
  BUFX2 U44 ( .A(n64), .Y(n46) );
  INVX1 U45 ( .A(n46), .Y(n78) );
  BUFX2 U46 ( .A(n65), .Y(n47) );
  INVX1 U47 ( .A(n47), .Y(n77) );
  BUFX2 U48 ( .A(n66), .Y(n48) );
  INVX1 U49 ( .A(n48), .Y(n76) );
  BUFX2 U50 ( .A(n67), .Y(n49) );
  INVX1 U51 ( .A(n49), .Y(n75) );
endmodule


module reg16_2 ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n1, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84;

  dff_47 d0 ( .q(\read<0> ), .d(n84), .clk(clk), .rst(rst) );
  dff_46 d1 ( .q(\read<1> ), .d(n83), .clk(clk), .rst(rst) );
  dff_45 d2 ( .q(\read<2> ), .d(n82), .clk(clk), .rst(rst) );
  dff_44 d3 ( .q(\read<3> ), .d(n81), .clk(clk), .rst(rst) );
  dff_43 d4 ( .q(\read<4> ), .d(n80), .clk(clk), .rst(rst) );
  dff_42 d5 ( .q(\read<5> ), .d(n79), .clk(clk), .rst(rst) );
  dff_41 d6 ( .q(\read<6> ), .d(n78), .clk(clk), .rst(rst) );
  dff_40 d7 ( .q(\read<7> ), .d(n77), .clk(clk), .rst(rst) );
  dff_39 d8 ( .q(\read<8> ), .d(n76), .clk(clk), .rst(rst) );
  dff_38 d9 ( .q(\read<9> ), .d(n75), .clk(clk), .rst(rst) );
  dff_37 d10 ( .q(\read<10> ), .d(n74), .clk(clk), .rst(rst) );
  dff_36 d11 ( .q(\read<11> ), .d(n73), .clk(clk), .rst(rst) );
  dff_35 d12 ( .q(\read<12> ), .d(n72), .clk(clk), .rst(rst) );
  dff_34 d13 ( .q(\read<13> ), .d(n71), .clk(clk), .rst(rst) );
  dff_33 d14 ( .q(\read<14> ), .d(n70), .clk(clk), .rst(rst) );
  dff_32 d15 ( .q(\read<15> ), .d(n69), .clk(clk), .rst(rst) );
  AOI22X1 U18 ( .A(\read<9> ), .B(n68), .C(\write<9> ), .D(n50), .Y(n67) );
  AOI22X1 U19 ( .A(\read<8> ), .B(n68), .C(\write<8> ), .D(n50), .Y(n66) );
  AOI22X1 U20 ( .A(\read<7> ), .B(n68), .C(\write<7> ), .D(n50), .Y(n65) );
  AOI22X1 U21 ( .A(\read<6> ), .B(n68), .C(\write<6> ), .D(n50), .Y(n64) );
  AOI22X1 U22 ( .A(\read<5> ), .B(n68), .C(\write<5> ), .D(n50), .Y(n63) );
  AOI22X1 U23 ( .A(\read<4> ), .B(n68), .C(\write<4> ), .D(n50), .Y(n62) );
  AOI22X1 U24 ( .A(\read<3> ), .B(n68), .C(\write<3> ), .D(n51), .Y(n61) );
  AOI22X1 U25 ( .A(\read<2> ), .B(n68), .C(\write<2> ), .D(n51), .Y(n60) );
  AOI22X1 U26 ( .A(\read<1> ), .B(n68), .C(\write<1> ), .D(n51), .Y(n59) );
  AOI22X1 U27 ( .A(\read<15> ), .B(n68), .C(\write<15> ), .D(n51), .Y(n58) );
  AOI22X1 U28 ( .A(\read<14> ), .B(n68), .C(\write<14> ), .D(n51), .Y(n57) );
  AOI22X1 U29 ( .A(\read<13> ), .B(n68), .C(\write<13> ), .D(n51), .Y(n56) );
  AOI22X1 U30 ( .A(\read<12> ), .B(n68), .C(\write<12> ), .D(n51), .Y(n55) );
  AOI22X1 U31 ( .A(\read<11> ), .B(n68), .C(\write<11> ), .D(n51), .Y(n54) );
  AOI22X1 U32 ( .A(\read<10> ), .B(n68), .C(\write<10> ), .D(n51), .Y(n53) );
  AOI22X1 U33 ( .A(\read<0> ), .B(n68), .C(\write<0> ), .D(n51), .Y(n52) );
  BUFX2 U1 ( .A(wr_en), .Y(n50) );
  BUFX2 U2 ( .A(wr_en), .Y(n51) );
  INVX1 U3 ( .A(n50), .Y(n68) );
  BUFX2 U4 ( .A(n52), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n84) );
  BUFX2 U6 ( .A(n53), .Y(n35) );
  INVX1 U7 ( .A(n35), .Y(n74) );
  BUFX2 U8 ( .A(n54), .Y(n36) );
  INVX1 U9 ( .A(n36), .Y(n73) );
  BUFX2 U10 ( .A(n55), .Y(n37) );
  INVX1 U11 ( .A(n37), .Y(n72) );
  BUFX2 U12 ( .A(n56), .Y(n38) );
  INVX1 U13 ( .A(n38), .Y(n71) );
  BUFX2 U14 ( .A(n57), .Y(n39) );
  INVX1 U15 ( .A(n39), .Y(n70) );
  BUFX2 U16 ( .A(n58), .Y(n40) );
  INVX1 U17 ( .A(n40), .Y(n69) );
  BUFX2 U34 ( .A(n59), .Y(n41) );
  INVX1 U35 ( .A(n41), .Y(n83) );
  BUFX2 U36 ( .A(n60), .Y(n42) );
  INVX1 U37 ( .A(n42), .Y(n82) );
  BUFX2 U38 ( .A(n61), .Y(n43) );
  INVX1 U39 ( .A(n43), .Y(n81) );
  BUFX2 U40 ( .A(n62), .Y(n44) );
  INVX1 U41 ( .A(n44), .Y(n80) );
  BUFX2 U42 ( .A(n63), .Y(n45) );
  INVX1 U43 ( .A(n45), .Y(n79) );
  BUFX2 U44 ( .A(n64), .Y(n46) );
  INVX1 U45 ( .A(n46), .Y(n78) );
  BUFX2 U46 ( .A(n65), .Y(n47) );
  INVX1 U47 ( .A(n47), .Y(n77) );
  BUFX2 U48 ( .A(n66), .Y(n48) );
  INVX1 U49 ( .A(n48), .Y(n76) );
  BUFX2 U50 ( .A(n67), .Y(n49) );
  INVX1 U51 ( .A(n49), .Y(n75) );
endmodule


module reg16_1 ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n1, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84;

  dff_31 d0 ( .q(\read<0> ), .d(n84), .clk(clk), .rst(rst) );
  dff_30 d1 ( .q(\read<1> ), .d(n83), .clk(clk), .rst(rst) );
  dff_29 d2 ( .q(\read<2> ), .d(n82), .clk(clk), .rst(rst) );
  dff_28 d3 ( .q(\read<3> ), .d(n81), .clk(clk), .rst(rst) );
  dff_27 d4 ( .q(\read<4> ), .d(n80), .clk(clk), .rst(rst) );
  dff_26 d5 ( .q(\read<5> ), .d(n79), .clk(clk), .rst(rst) );
  dff_25 d6 ( .q(\read<6> ), .d(n78), .clk(clk), .rst(rst) );
  dff_24 d7 ( .q(\read<7> ), .d(n77), .clk(clk), .rst(rst) );
  dff_23 d8 ( .q(\read<8> ), .d(n76), .clk(clk), .rst(rst) );
  dff_22 d9 ( .q(\read<9> ), .d(n75), .clk(clk), .rst(rst) );
  dff_21 d10 ( .q(\read<10> ), .d(n74), .clk(clk), .rst(rst) );
  dff_20 d11 ( .q(\read<11> ), .d(n73), .clk(clk), .rst(rst) );
  dff_19 d12 ( .q(\read<12> ), .d(n72), .clk(clk), .rst(rst) );
  dff_18 d13 ( .q(\read<13> ), .d(n71), .clk(clk), .rst(rst) );
  dff_17 d14 ( .q(\read<14> ), .d(n70), .clk(clk), .rst(rst) );
  dff_16 d15 ( .q(\read<15> ), .d(n69), .clk(clk), .rst(rst) );
  AOI22X1 U18 ( .A(\read<9> ), .B(n68), .C(\write<9> ), .D(n50), .Y(n67) );
  AOI22X1 U19 ( .A(\read<8> ), .B(n68), .C(\write<8> ), .D(n50), .Y(n66) );
  AOI22X1 U20 ( .A(\read<7> ), .B(n68), .C(\write<7> ), .D(n50), .Y(n65) );
  AOI22X1 U21 ( .A(\read<6> ), .B(n68), .C(\write<6> ), .D(n50), .Y(n64) );
  AOI22X1 U22 ( .A(\read<5> ), .B(n68), .C(\write<5> ), .D(n50), .Y(n63) );
  AOI22X1 U23 ( .A(\read<4> ), .B(n68), .C(\write<4> ), .D(n50), .Y(n62) );
  AOI22X1 U24 ( .A(\read<3> ), .B(n68), .C(\write<3> ), .D(n51), .Y(n61) );
  AOI22X1 U25 ( .A(\read<2> ), .B(n68), .C(\write<2> ), .D(n51), .Y(n60) );
  AOI22X1 U26 ( .A(\read<1> ), .B(n68), .C(\write<1> ), .D(n51), .Y(n59) );
  AOI22X1 U27 ( .A(\read<15> ), .B(n68), .C(\write<15> ), .D(n51), .Y(n58) );
  AOI22X1 U28 ( .A(\read<14> ), .B(n68), .C(\write<14> ), .D(n51), .Y(n57) );
  AOI22X1 U29 ( .A(\read<13> ), .B(n68), .C(\write<13> ), .D(n51), .Y(n56) );
  AOI22X1 U30 ( .A(\read<12> ), .B(n68), .C(\write<12> ), .D(n51), .Y(n55) );
  AOI22X1 U31 ( .A(\read<11> ), .B(n68), .C(\write<11> ), .D(n51), .Y(n54) );
  AOI22X1 U32 ( .A(\read<10> ), .B(n68), .C(\write<10> ), .D(n51), .Y(n53) );
  AOI22X1 U33 ( .A(\read<0> ), .B(n68), .C(\write<0> ), .D(n51), .Y(n52) );
  BUFX2 U1 ( .A(wr_en), .Y(n50) );
  BUFX2 U2 ( .A(wr_en), .Y(n51) );
  INVX1 U3 ( .A(n50), .Y(n68) );
  BUFX2 U4 ( .A(n52), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n84) );
  BUFX2 U6 ( .A(n53), .Y(n35) );
  INVX1 U7 ( .A(n35), .Y(n74) );
  BUFX2 U8 ( .A(n54), .Y(n36) );
  INVX1 U9 ( .A(n36), .Y(n73) );
  BUFX2 U10 ( .A(n55), .Y(n37) );
  INVX1 U11 ( .A(n37), .Y(n72) );
  BUFX2 U12 ( .A(n56), .Y(n38) );
  INVX1 U13 ( .A(n38), .Y(n71) );
  BUFX2 U14 ( .A(n57), .Y(n39) );
  INVX1 U15 ( .A(n39), .Y(n70) );
  BUFX2 U16 ( .A(n58), .Y(n40) );
  INVX1 U17 ( .A(n40), .Y(n69) );
  BUFX2 U34 ( .A(n59), .Y(n41) );
  INVX1 U35 ( .A(n41), .Y(n83) );
  BUFX2 U36 ( .A(n60), .Y(n42) );
  INVX1 U37 ( .A(n42), .Y(n82) );
  BUFX2 U38 ( .A(n61), .Y(n43) );
  INVX1 U39 ( .A(n43), .Y(n81) );
  BUFX2 U40 ( .A(n62), .Y(n44) );
  INVX1 U41 ( .A(n44), .Y(n80) );
  BUFX2 U42 ( .A(n63), .Y(n45) );
  INVX1 U43 ( .A(n45), .Y(n79) );
  BUFX2 U44 ( .A(n64), .Y(n46) );
  INVX1 U45 ( .A(n46), .Y(n78) );
  BUFX2 U46 ( .A(n65), .Y(n47) );
  INVX1 U47 ( .A(n47), .Y(n77) );
  BUFX2 U48 ( .A(n66), .Y(n48) );
  INVX1 U49 ( .A(n48), .Y(n76) );
  BUFX2 U50 ( .A(n67), .Y(n49) );
  INVX1 U51 ( .A(n49), .Y(n75) );
endmodule


module reg16_0 ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n1, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84;

  dff_15 d0 ( .q(\read<0> ), .d(n84), .clk(clk), .rst(rst) );
  dff_14 d1 ( .q(\read<1> ), .d(n83), .clk(clk), .rst(rst) );
  dff_13 d2 ( .q(\read<2> ), .d(n82), .clk(clk), .rst(rst) );
  dff_12 d3 ( .q(\read<3> ), .d(n81), .clk(clk), .rst(rst) );
  dff_11 d4 ( .q(\read<4> ), .d(n80), .clk(clk), .rst(rst) );
  dff_10 d5 ( .q(\read<5> ), .d(n79), .clk(clk), .rst(rst) );
  dff_9 d6 ( .q(\read<6> ), .d(n78), .clk(clk), .rst(rst) );
  dff_8 d7 ( .q(\read<7> ), .d(n77), .clk(clk), .rst(rst) );
  dff_7 d8 ( .q(\read<8> ), .d(n76), .clk(clk), .rst(rst) );
  dff_6 d9 ( .q(\read<9> ), .d(n75), .clk(clk), .rst(rst) );
  dff_5 d10 ( .q(\read<10> ), .d(n74), .clk(clk), .rst(rst) );
  dff_4 d11 ( .q(\read<11> ), .d(n73), .clk(clk), .rst(rst) );
  dff_3 d12 ( .q(\read<12> ), .d(n72), .clk(clk), .rst(rst) );
  dff_2 d13 ( .q(\read<13> ), .d(n71), .clk(clk), .rst(rst) );
  dff_1 d14 ( .q(\read<14> ), .d(n70), .clk(clk), .rst(rst) );
  dff_0 d15 ( .q(\read<15> ), .d(n69), .clk(clk), .rst(rst) );
  AOI22X1 U18 ( .A(\read<9> ), .B(n68), .C(\write<9> ), .D(n50), .Y(n67) );
  AOI22X1 U19 ( .A(\read<8> ), .B(n68), .C(\write<8> ), .D(n50), .Y(n66) );
  AOI22X1 U20 ( .A(\read<7> ), .B(n68), .C(\write<7> ), .D(n50), .Y(n65) );
  AOI22X1 U21 ( .A(\read<6> ), .B(n68), .C(\write<6> ), .D(n50), .Y(n64) );
  AOI22X1 U22 ( .A(\read<5> ), .B(n68), .C(\write<5> ), .D(n50), .Y(n63) );
  AOI22X1 U23 ( .A(\read<4> ), .B(n68), .C(\write<4> ), .D(n50), .Y(n62) );
  AOI22X1 U24 ( .A(\read<3> ), .B(n68), .C(\write<3> ), .D(n51), .Y(n61) );
  AOI22X1 U25 ( .A(\read<2> ), .B(n68), .C(\write<2> ), .D(n51), .Y(n60) );
  AOI22X1 U26 ( .A(\read<1> ), .B(n68), .C(\write<1> ), .D(n51), .Y(n59) );
  AOI22X1 U27 ( .A(\read<15> ), .B(n68), .C(\write<15> ), .D(n51), .Y(n58) );
  AOI22X1 U28 ( .A(\read<14> ), .B(n68), .C(\write<14> ), .D(n51), .Y(n57) );
  AOI22X1 U29 ( .A(\read<13> ), .B(n68), .C(\write<13> ), .D(n51), .Y(n56) );
  AOI22X1 U30 ( .A(\read<12> ), .B(n68), .C(\write<12> ), .D(n51), .Y(n55) );
  AOI22X1 U31 ( .A(\read<11> ), .B(n68), .C(\write<11> ), .D(n51), .Y(n54) );
  AOI22X1 U32 ( .A(\read<10> ), .B(n68), .C(\write<10> ), .D(n51), .Y(n53) );
  AOI22X1 U33 ( .A(\read<0> ), .B(n68), .C(\write<0> ), .D(n51), .Y(n52) );
  BUFX2 U1 ( .A(wr_en), .Y(n50) );
  BUFX2 U2 ( .A(wr_en), .Y(n51) );
  INVX1 U3 ( .A(n50), .Y(n68) );
  BUFX2 U4 ( .A(n52), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n84) );
  BUFX2 U6 ( .A(n53), .Y(n35) );
  INVX1 U7 ( .A(n35), .Y(n74) );
  BUFX2 U8 ( .A(n54), .Y(n36) );
  INVX1 U9 ( .A(n36), .Y(n73) );
  BUFX2 U10 ( .A(n55), .Y(n37) );
  INVX1 U11 ( .A(n37), .Y(n72) );
  BUFX2 U12 ( .A(n56), .Y(n38) );
  INVX1 U13 ( .A(n38), .Y(n71) );
  BUFX2 U14 ( .A(n57), .Y(n39) );
  INVX1 U15 ( .A(n39), .Y(n70) );
  BUFX2 U16 ( .A(n58), .Y(n40) );
  INVX1 U17 ( .A(n40), .Y(n69) );
  BUFX2 U34 ( .A(n59), .Y(n41) );
  INVX1 U35 ( .A(n41), .Y(n83) );
  BUFX2 U36 ( .A(n60), .Y(n42) );
  INVX1 U37 ( .A(n42), .Y(n82) );
  BUFX2 U38 ( .A(n61), .Y(n43) );
  INVX1 U39 ( .A(n43), .Y(n81) );
  BUFX2 U40 ( .A(n62), .Y(n44) );
  INVX1 U41 ( .A(n44), .Y(n80) );
  BUFX2 U42 ( .A(n63), .Y(n45) );
  INVX1 U43 ( .A(n45), .Y(n79) );
  BUFX2 U44 ( .A(n64), .Y(n46) );
  INVX1 U45 ( .A(n46), .Y(n78) );
  BUFX2 U46 ( .A(n65), .Y(n47) );
  INVX1 U47 ( .A(n47), .Y(n77) );
  BUFX2 U48 ( .A(n66), .Y(n48) );
  INVX1 U49 ( .A(n48), .Y(n76) );
  BUFX2 U50 ( .A(n67), .Y(n49) );
  INVX1 U51 ( .A(n49), .Y(n75) );
endmodule


module CLA4_3 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, Cout, P, G, .S({\S<3> , \S<2> , \S<1> , \S<0> }
        ) );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output Cout, P, G, \S<3> , \S<2> , \S<1> , \S<0> ;
  wire   p0, g0, p1, g1, p2, g2, c3, p3, g3, n1, n2, n3, n4, n5, n6, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42;

  pfa_15 bit0 ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(p0), .G(g0)
         );
  pfa_14 bit1 ( .A(\A<1> ), .B(\B<1> ), .Cin(n20), .S(\S<1> ), .P(p1), .G(g1)
         );
  pfa_13 bit2 ( .A(\A<2> ), .B(\B<2> ), .Cin(n42), .S(\S<2> ), .P(p2), .G(g2)
         );
  pfa_12 bit3 ( .A(\A<3> ), .B(\B<3> ), .Cin(c3), .S(\S<3> ), .P(p3), .G(g3)
         );
  INVX2 U1 ( .A(p2), .Y(n36) );
  INVX1 U2 ( .A(n31), .Y(n1) );
  INVX1 U3 ( .A(g0), .Y(n34) );
  INVX1 U4 ( .A(Cin), .Y(n40) );
  INVX1 U5 ( .A(g3), .Y(n2) );
  INVX1 U6 ( .A(n2), .Y(n3) );
  AND2X2 U7 ( .A(n1), .B(Cin), .Y(n11) );
  BUFX2 U8 ( .A(P), .Y(n4) );
  BUFX2 U9 ( .A(G), .Y(n5) );
  INVX1 U10 ( .A(n6), .Y(n37) );
  NOR3X1 U11 ( .A(n3), .B(n14), .C(n25), .Y(n6) );
  AND2X2 U12 ( .A(n37), .B(n22), .Y(G) );
  INVX1 U13 ( .A(g2), .Y(n8) );
  OR2X2 U14 ( .A(g1), .B(n27), .Y(n24) );
  INVX1 U15 ( .A(g1), .Y(n33) );
  AND2X2 U16 ( .A(p1), .B(g0), .Y(n25) );
  AND2X2 U17 ( .A(p2), .B(p3), .Y(n9) );
  INVX1 U18 ( .A(n9), .Y(n10) );
  INVX1 U19 ( .A(n11), .Y(n12) );
  OR2X2 U20 ( .A(p3), .B(g3), .Y(n13) );
  OR2X2 U21 ( .A(g2), .B(g1), .Y(n14) );
  BUFX2 U22 ( .A(n35), .Y(n15) );
  OR2X2 U23 ( .A(g2), .B(g3), .Y(n16) );
  INVX1 U24 ( .A(n16), .Y(n17) );
  BUFX2 U25 ( .A(n32), .Y(n18) );
  AND2X2 U26 ( .A(n34), .B(n12), .Y(n19) );
  INVX1 U27 ( .A(n19), .Y(n20) );
  INVX1 U28 ( .A(n38), .Y(n21) );
  INVX1 U29 ( .A(n21), .Y(n22) );
  INVX1 U30 ( .A(n13), .Y(n23) );
  INVX1 U31 ( .A(n11), .Y(n26) );
  INVX1 U32 ( .A(n5), .Y(n39) );
  INVX1 U33 ( .A(n30), .Y(n27) );
  INVX1 U34 ( .A(p0), .Y(n31) );
  BUFX2 U35 ( .A(n36), .Y(n28) );
  INVX1 U36 ( .A(p1), .Y(n30) );
  NOR3X1 U37 ( .A(n30), .B(n31), .C(n10), .Y(P) );
  INVX1 U38 ( .A(n4), .Y(n41) );
  AOI21X1 U39 ( .A(n27), .B(n20), .C(g1), .Y(n32) );
  OAI21X1 U40 ( .A(n18), .B(n28), .C(n8), .Y(c3) );
  NAND3X1 U41 ( .A(n34), .B(n26), .C(n33), .Y(n35) );
  AND2X2 U42 ( .A(n15), .B(n24), .Y(n42) );
  AOI21X1 U43 ( .A(n36), .B(n17), .C(n23), .Y(n38) );
  OAI21X1 U44 ( .A(n41), .B(n40), .C(n39), .Y(Cout) );
endmodule


module CLA4_2 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, Cout, P, G, .S({\S<3> , \S<2> , \S<1> , \S<0> }
        ) );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output Cout, P, G, \S<3> , \S<2> , \S<1> , \S<0> ;
  wire   p0, g0, p1, g1, p2, g2, p3, g3, n1, n2, n3, n4, n5, n6, n7, n8, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51;

  pfa_11 bit0 ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(p0), .G(g0)
         );
  pfa_10 bit1 ( .A(\A<1> ), .B(\B<1> ), .Cin(n50), .S(\S<1> ), .P(p1), .G(g1)
         );
  pfa_9 bit2 ( .A(\A<2> ), .B(\B<2> ), .Cin(n48), .S(\S<2> ), .P(p2), .G(g2)
         );
  pfa_8 bit3 ( .A(\A<3> ), .B(\B<3> ), .Cin(n49), .S(\S<3> ), .P(p3), .G(g3)
         );
  INVX1 U1 ( .A(p3), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(n2) );
  INVX1 U3 ( .A(g0), .Y(n34) );
  INVX1 U4 ( .A(g2), .Y(n42) );
  INVX1 U5 ( .A(n34), .Y(n12) );
  INVX1 U6 ( .A(n26), .Y(n3) );
  AND2X2 U7 ( .A(n38), .B(n34), .Y(n4) );
  BUFX2 U8 ( .A(p1), .Y(n5) );
  INVX1 U9 ( .A(n43), .Y(n6) );
  INVX1 U10 ( .A(n47), .Y(n7) );
  AND2X2 U11 ( .A(Cin), .B(n30), .Y(n26) );
  INVX1 U12 ( .A(g3), .Y(n47) );
  AND2X2 U13 ( .A(n27), .B(n4), .Y(n15) );
  BUFX2 U14 ( .A(Cin), .Y(n8) );
  INVX1 U15 ( .A(g1), .Y(n38) );
  AND2X2 U16 ( .A(n10), .B(p0), .Y(P) );
  INVX1 U17 ( .A(n40), .Y(n10) );
  AND2X2 U18 ( .A(n6), .B(p1), .Y(n23) );
  OAI21X1 U19 ( .A(n30), .B(n12), .C(n19), .Y(n11) );
  INVX1 U20 ( .A(n11), .Y(n50) );
  AND2X2 U21 ( .A(n36), .B(n43), .Y(n13) );
  INVX1 U22 ( .A(n13), .Y(n14) );
  INVX1 U23 ( .A(n15), .Y(n16) );
  INVX1 U24 ( .A(p2), .Y(n43) );
  BUFX2 U25 ( .A(n31), .Y(n17) );
  INVX1 U26 ( .A(n35), .Y(n36) );
  BUFX2 U27 ( .A(n46), .Y(n18) );
  OR2X2 U28 ( .A(Cin), .B(g0), .Y(n19) );
  INVX1 U29 ( .A(n39), .Y(n20) );
  INVX1 U30 ( .A(n20), .Y(n21) );
  BUFX2 U31 ( .A(n44), .Y(n22) );
  INVX1 U32 ( .A(n23), .Y(n24) );
  BUFX2 U33 ( .A(P), .Y(n25) );
  INVX1 U34 ( .A(n26), .Y(n27) );
  INVX1 U35 ( .A(n51), .Y(n28) );
  INVX1 U36 ( .A(n28), .Y(G) );
  INVX1 U37 ( .A(p0), .Y(n41) );
  INVX1 U38 ( .A(n41), .Y(n30) );
  AND2X2 U39 ( .A(n3), .B(n34), .Y(n32) );
  AOI21X1 U40 ( .A(g1), .B(n6), .C(g2), .Y(n31) );
  OAI21X1 U41 ( .A(n32), .B(n24), .C(n17), .Y(n49) );
  OR2X2 U42 ( .A(p1), .B(g1), .Y(n33) );
  AND2X2 U43 ( .A(n16), .B(n33), .Y(n48) );
  OR2X2 U44 ( .A(g3), .B(g2), .Y(n35) );
  AOI21X1 U45 ( .A(g0), .B(p1), .C(n35), .Y(n39) );
  OAI21X1 U46 ( .A(n7), .B(n2), .C(n14), .Y(n37) );
  AOI21X1 U47 ( .A(n38), .B(n21), .C(n37), .Y(n51) );
  NAND3X1 U48 ( .A(p1), .B(p2), .C(p3), .Y(n40) );
  AOI21X1 U49 ( .A(n12), .B(n5), .C(g1), .Y(n44) );
  OAI21X1 U50 ( .A(n22), .B(n43), .C(n42), .Y(n45) );
  AOI22X1 U51 ( .A(n2), .B(n45), .C(n25), .D(n8), .Y(n46) );
  NAND2X1 U52 ( .A(n47), .B(n18), .Y(Cout) );
endmodule


module CLA4_1 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, Cout, P, G, .S({\S<3> , \S<2> , \S<1> , \S<0> }
        ) );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output Cout, P, G, \S<3> , \S<2> , \S<1> , \S<0> ;
  wire   p0, g0, p1, g1, p2, g2, c3, p3, g3, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58;

  pfa_7 bit0 ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(p0), .G(g0)
         );
  pfa_6 bit1 ( .A(\A<1> ), .B(\B<1> ), .Cin(n28), .S(\S<1> ), .P(p1), .G(g1)
         );
  pfa_5 bit2 ( .A(\A<2> ), .B(\B<2> ), .Cin(n39), .S(\S<2> ), .P(p2), .G(g2)
         );
  pfa_4 bit3 ( .A(\A<3> ), .B(\B<3> ), .Cin(n40), .S(\S<3> ), .P(p3), .G(g3)
         );
  BUFX2 U1 ( .A(g1), .Y(n1) );
  INVX1 U2 ( .A(p0), .Y(n2) );
  INVX1 U3 ( .A(n2), .Y(n3) );
  INVX1 U4 ( .A(n55), .Y(n4) );
  BUFX2 U5 ( .A(Cin), .Y(n5) );
  BUFX2 U6 ( .A(p1), .Y(n6) );
  OR2X2 U7 ( .A(n3), .B(g0), .Y(n34) );
  AND2X2 U8 ( .A(n6), .B(n3), .Y(n43) );
  AND2X2 U9 ( .A(g0), .B(n6), .Y(n18) );
  OR2X2 U10 ( .A(Cin), .B(g0), .Y(n25) );
  OR2X2 U11 ( .A(n35), .B(n26), .Y(n27) );
  OR2X2 U12 ( .A(n52), .B(n51), .Y(n11) );
  AND2X2 U13 ( .A(Cin), .B(n21), .Y(n22) );
  OR2X2 U14 ( .A(g1), .B(g3), .Y(n10) );
  NOR3X1 U15 ( .A(n4), .B(p1), .C(n10), .Y(n7) );
  INVX1 U16 ( .A(g2), .Y(n55) );
  OR2X2 U17 ( .A(Cin), .B(n46), .Y(n24) );
  OR2X2 U18 ( .A(g1), .B(g2), .Y(n12) );
  OR2X2 U19 ( .A(g2), .B(g3), .Y(n8) );
  INVX1 U20 ( .A(n8), .Y(n9) );
  INVX1 U21 ( .A(n12), .Y(n13) );
  BUFX2 U22 ( .A(n53), .Y(n14) );
  OR2X2 U23 ( .A(n14), .B(n54), .Y(n15) );
  INVX1 U24 ( .A(n15), .Y(P) );
  INVX1 U25 ( .A(n15), .Y(n17) );
  INVX1 U26 ( .A(n18), .Y(n19) );
  INVX1 U27 ( .A(n7), .Y(n20) );
  AND2X1 U28 ( .A(p2), .B(n43), .Y(n21) );
  INVX1 U29 ( .A(n22), .Y(n23) );
  INVX1 U30 ( .A(n25), .Y(n26) );
  INVX1 U31 ( .A(n27), .Y(n28) );
  AND2X2 U32 ( .A(n13), .B(n57), .Y(n29) );
  INVX1 U33 ( .A(n29), .Y(n30) );
  AND2X2 U34 ( .A(n50), .B(n9), .Y(n31) );
  INVX1 U35 ( .A(n31), .Y(n32) );
  BUFX2 U36 ( .A(n56), .Y(n33) );
  INVX1 U37 ( .A(n34), .Y(n35) );
  INVX1 U38 ( .A(n24), .Y(n36) );
  AND2X1 U39 ( .A(n55), .B(n45), .Y(n37) );
  INVX1 U40 ( .A(n37), .Y(n38) );
  BUFX2 U41 ( .A(n58), .Y(n39) );
  BUFX2 U42 ( .A(c3), .Y(n40) );
  INVX1 U43 ( .A(n11), .Y(G) );
  INVX1 U44 ( .A(n43), .Y(n42) );
  AND2X1 U45 ( .A(p2), .B(n46), .Y(n44) );
  INVX1 U46 ( .A(n44), .Y(n45) );
  INVX1 U47 ( .A(n47), .Y(n46) );
  AND2X2 U48 ( .A(n49), .B(n19), .Y(n47) );
  INVX1 U49 ( .A(p2), .Y(n50) );
  INVX1 U50 ( .A(n1), .Y(n49) );
  INVX1 U51 ( .A(n6), .Y(n54) );
  INVX1 U52 ( .A(n57), .Y(n48) );
  INVX1 U53 ( .A(g3), .Y(n57) );
  NAND3X1 U54 ( .A(n55), .B(n45), .C(n23), .Y(c3) );
  AOI21X1 U55 ( .A(n42), .B(n47), .C(n36), .Y(n58) );
  OAI21X1 U56 ( .A(g0), .B(n30), .C(n32), .Y(n52) );
  OAI21X1 U57 ( .A(n48), .B(p3), .C(n20), .Y(n51) );
  NAND3X1 U58 ( .A(p3), .B(p2), .C(p0), .Y(n53) );
  AOI22X1 U59 ( .A(p3), .B(n38), .C(n5), .D(n17), .Y(n56) );
  NAND2X1 U60 ( .A(n57), .B(n33), .Y(Cout) );
endmodule


module CLA4_0 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, Cout, P, G, .S({\S<3> , \S<2> , \S<1> , \S<0> }
        ) );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output Cout, P, G, \S<3> , \S<2> , \S<1> , \S<0> ;
  wire   p0, g0, p1, g1, p2, g2, p3, g3, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46;

  pfa_3 bit0 ( .A(\A<0> ), .B(\B<0> ), .Cin(n35), .S(\S<0> ), .P(p0), .G(g0)
         );
  pfa_2 bit1 ( .A(\A<1> ), .B(\B<1> ), .Cin(n11), .S(\S<1> ), .P(p1), .G(g1)
         );
  pfa_1 bit2 ( .A(\A<2> ), .B(\B<2> ), .Cin(n28), .S(\S<2> ), .P(p2), .G(g2)
         );
  pfa_0 bit3 ( .A(\A<3> ), .B(\B<3> ), .Cin(n13), .S(\S<3> ), .P(p3), .G(g3)
         );
  INVX2 U1 ( .A(n37), .Y(n40) );
  INVX1 U2 ( .A(n36), .Y(n39) );
  INVX1 U3 ( .A(g2), .Y(n42) );
  INVX1 U4 ( .A(g3), .Y(n45) );
  BUFX2 U5 ( .A(p2), .Y(n1) );
  INVX1 U6 ( .A(n34), .Y(n2) );
  OAI21X1 U7 ( .A(n39), .B(n38), .C(n37), .Y(n3) );
  AND2X2 U8 ( .A(p0), .B(n3), .Y(n20) );
  INVX1 U9 ( .A(n34), .Y(n35) );
  AND2X2 U10 ( .A(n33), .B(n21), .Y(n12) );
  AND2X2 U11 ( .A(n2), .B(P), .Y(n22) );
  AND2X2 U12 ( .A(n2), .B(n26), .Y(n14) );
  OR2X2 U13 ( .A(n2), .B(g0), .Y(n8) );
  AND2X2 U14 ( .A(p3), .B(n44), .Y(n4) );
  INVX1 U15 ( .A(n4), .Y(n5) );
  AND2X2 U16 ( .A(n41), .B(n34), .Y(n6) );
  INVX1 U17 ( .A(n6), .Y(n7) );
  INVX1 U18 ( .A(n8), .Y(n9) );
  OR2X2 U19 ( .A(n9), .B(n25), .Y(n10) );
  INVX1 U20 ( .A(n10), .Y(n11) );
  AND2X2 U21 ( .A(n7), .B(n19), .Y(n13) );
  INVX1 U22 ( .A(n14), .Y(n15) );
  INVX1 U23 ( .A(n18), .Y(n16) );
  INVX1 U24 ( .A(n16), .Y(n17) );
  BUFX2 U25 ( .A(n29), .Y(n18) );
  INVX1 U26 ( .A(n12), .Y(n19) );
  INVX1 U27 ( .A(n20), .Y(n21) );
  INVX1 U28 ( .A(n22), .Y(n23) );
  OR2X1 U29 ( .A(g0), .B(p0), .Y(n24) );
  INVX1 U30 ( .A(n24), .Y(n25) );
  INVX1 U31 ( .A(n46), .Y(P) );
  AND2X1 U32 ( .A(p0), .B(p1), .Y(n26) );
  AND2X2 U33 ( .A(n15), .B(n17), .Y(n27) );
  INVX1 U34 ( .A(n27), .Y(n28) );
  AOI21X1 U35 ( .A(g0), .B(p1), .C(g1), .Y(n29) );
  AND2X2 U36 ( .A(n45), .B(n5), .Y(n30) );
  INVX1 U37 ( .A(n30), .Y(G) );
  INVX1 U38 ( .A(n41), .Y(n32) );
  INVX1 U39 ( .A(n32), .Y(n33) );
  INVX1 U40 ( .A(n1), .Y(n43) );
  INVX1 U41 ( .A(p1), .Y(n38) );
  INVX1 U42 ( .A(Cin), .Y(n34) );
  OR2X2 U43 ( .A(p2), .B(g2), .Y(n36) );
  OAI21X1 U44 ( .A(g2), .B(g1), .C(n36), .Y(n37) );
  OAI21X1 U45 ( .A(g0), .B(n40), .C(n3), .Y(n41) );
  OAI21X1 U46 ( .A(n18), .B(n43), .C(n42), .Y(n44) );
  NAND3X1 U47 ( .A(p3), .B(n1), .C(n26), .Y(n46) );
  NAND2X1 U48 ( .A(n30), .B(n23), .Y(Cout) );
endmodule


module dff_664 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_663 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_662 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_661 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_660 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_659 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_658 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_657 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_656 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_655 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_654 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_653 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_652 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_651 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_650 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_649 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_648 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module reg16_9 ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n1, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85;

  dff_159 d0 ( .q(\read<0> ), .d(n85), .clk(clk), .rst(rst) );
  dff_158 d1 ( .q(\read<1> ), .d(n84), .clk(clk), .rst(rst) );
  dff_157 d2 ( .q(\read<2> ), .d(n83), .clk(clk), .rst(rst) );
  dff_156 d3 ( .q(\read<3> ), .d(n82), .clk(clk), .rst(rst) );
  dff_155 d4 ( .q(\read<4> ), .d(n81), .clk(clk), .rst(rst) );
  dff_154 d5 ( .q(\read<5> ), .d(n80), .clk(clk), .rst(rst) );
  dff_153 d6 ( .q(\read<6> ), .d(n79), .clk(clk), .rst(rst) );
  dff_152 d7 ( .q(\read<7> ), .d(n78), .clk(clk), .rst(rst) );
  dff_151 d8 ( .q(\read<8> ), .d(n77), .clk(clk), .rst(rst) );
  dff_150 d9 ( .q(\read<9> ), .d(n76), .clk(clk), .rst(rst) );
  dff_149 d10 ( .q(\read<10> ), .d(n75), .clk(clk), .rst(rst) );
  dff_148 d11 ( .q(\read<11> ), .d(n74), .clk(clk), .rst(rst) );
  dff_147 d12 ( .q(\read<12> ), .d(n73), .clk(clk), .rst(rst) );
  dff_146 d13 ( .q(\read<13> ), .d(n72), .clk(clk), .rst(rst) );
  dff_145 d14 ( .q(\read<14> ), .d(n71), .clk(clk), .rst(rst) );
  dff_144 d15 ( .q(\read<15> ), .d(n70), .clk(clk), .rst(rst) );
  AOI22X1 U18 ( .A(\read<9> ), .B(n69), .C(\write<9> ), .D(n51), .Y(n68) );
  AOI22X1 U19 ( .A(\read<8> ), .B(n69), .C(\write<8> ), .D(n51), .Y(n67) );
  AOI22X1 U20 ( .A(\read<7> ), .B(n69), .C(\write<7> ), .D(n51), .Y(n66) );
  AOI22X1 U21 ( .A(\read<6> ), .B(n69), .C(\write<6> ), .D(n51), .Y(n65) );
  AOI22X1 U22 ( .A(\read<5> ), .B(n69), .C(\write<5> ), .D(n51), .Y(n64) );
  AOI22X1 U23 ( .A(\read<4> ), .B(n69), .C(\write<4> ), .D(n51), .Y(n63) );
  AOI22X1 U24 ( .A(\read<3> ), .B(n69), .C(\write<3> ), .D(n52), .Y(n62) );
  AOI22X1 U25 ( .A(\read<2> ), .B(n69), .C(\write<2> ), .D(n52), .Y(n61) );
  AOI22X1 U26 ( .A(n1), .B(n69), .C(\write<1> ), .D(n52), .Y(n60) );
  AOI22X1 U27 ( .A(\read<15> ), .B(n69), .C(\write<15> ), .D(n52), .Y(n59) );
  AOI22X1 U28 ( .A(\read<14> ), .B(n69), .C(\write<14> ), .D(n52), .Y(n58) );
  AOI22X1 U29 ( .A(\read<13> ), .B(n69), .C(\write<13> ), .D(n52), .Y(n57) );
  AOI22X1 U30 ( .A(\read<12> ), .B(n69), .C(\write<12> ), .D(n52), .Y(n56) );
  AOI22X1 U31 ( .A(\read<11> ), .B(n69), .C(\write<11> ), .D(n52), .Y(n55) );
  AOI22X1 U32 ( .A(\read<10> ), .B(n69), .C(\write<10> ), .D(n52), .Y(n54) );
  AOI22X1 U33 ( .A(\read<0> ), .B(n69), .C(\write<0> ), .D(n52), .Y(n53) );
  BUFX2 U1 ( .A(wr_en), .Y(n51) );
  BUFX2 U2 ( .A(wr_en), .Y(n52) );
  BUFX2 U3 ( .A(\read<1> ), .Y(n1) );
  INVX1 U4 ( .A(n51), .Y(n69) );
  BUFX2 U5 ( .A(n53), .Y(n35) );
  INVX1 U6 ( .A(n35), .Y(n85) );
  BUFX2 U7 ( .A(n54), .Y(n36) );
  INVX1 U8 ( .A(n36), .Y(n75) );
  BUFX2 U9 ( .A(n55), .Y(n37) );
  INVX1 U10 ( .A(n37), .Y(n74) );
  BUFX2 U11 ( .A(n56), .Y(n38) );
  INVX1 U12 ( .A(n38), .Y(n73) );
  BUFX2 U13 ( .A(n57), .Y(n39) );
  INVX1 U14 ( .A(n39), .Y(n72) );
  BUFX2 U15 ( .A(n58), .Y(n40) );
  INVX1 U16 ( .A(n40), .Y(n71) );
  BUFX2 U17 ( .A(n59), .Y(n41) );
  INVX1 U34 ( .A(n41), .Y(n70) );
  BUFX2 U35 ( .A(n60), .Y(n42) );
  INVX1 U36 ( .A(n42), .Y(n84) );
  BUFX2 U37 ( .A(n61), .Y(n43) );
  INVX1 U38 ( .A(n43), .Y(n83) );
  BUFX2 U39 ( .A(n62), .Y(n44) );
  INVX1 U40 ( .A(n44), .Y(n82) );
  BUFX2 U41 ( .A(n63), .Y(n45) );
  INVX1 U42 ( .A(n45), .Y(n81) );
  BUFX2 U43 ( .A(n64), .Y(n46) );
  INVX1 U44 ( .A(n46), .Y(n80) );
  BUFX2 U45 ( .A(n65), .Y(n47) );
  INVX1 U46 ( .A(n47), .Y(n79) );
  BUFX2 U47 ( .A(n66), .Y(n48) );
  INVX1 U48 ( .A(n48), .Y(n78) );
  BUFX2 U49 ( .A(n67), .Y(n49) );
  INVX1 U50 ( .A(n49), .Y(n77) );
  BUFX2 U51 ( .A(n68), .Y(n50) );
  INVX1 U52 ( .A(n50), .Y(n76) );
endmodule


module reg16_8 ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54;

  dff_143 d0 ( .q(\read<0> ), .d(n39), .clk(clk), .rst(rst) );
  dff_142 d1 ( .q(\read<1> ), .d(n40), .clk(clk), .rst(rst) );
  dff_141 d2 ( .q(\read<2> ), .d(n41), .clk(clk), .rst(rst) );
  dff_140 d3 ( .q(\read<3> ), .d(n42), .clk(clk), .rst(rst) );
  dff_139 d4 ( .q(\read<4> ), .d(n43), .clk(clk), .rst(rst) );
  dff_138 d5 ( .q(\read<5> ), .d(n44), .clk(clk), .rst(rst) );
  dff_137 d6 ( .q(\read<6> ), .d(n45), .clk(clk), .rst(rst) );
  dff_136 d7 ( .q(\read<7> ), .d(n46), .clk(clk), .rst(rst) );
  dff_135 d8 ( .q(\read<8> ), .d(n47), .clk(clk), .rst(rst) );
  dff_134 d9 ( .q(\read<9> ), .d(n48), .clk(clk), .rst(rst) );
  dff_133 d10 ( .q(\read<10> ), .d(n49), .clk(clk), .rst(rst) );
  dff_132 d11 ( .q(\read<11> ), .d(n50), .clk(clk), .rst(rst) );
  dff_131 d12 ( .q(\read<12> ), .d(n51), .clk(clk), .rst(rst) );
  dff_130 d13 ( .q(\read<13> ), .d(n52), .clk(clk), .rst(rst) );
  dff_129 d14 ( .q(\read<14> ), .d(n53), .clk(clk), .rst(rst) );
  dff_128 d15 ( .q(\read<15> ), .d(n54), .clk(clk), .rst(rst) );
  INVX1 U1 ( .A(\read<6> ), .Y(n26) );
  INVX1 U2 ( .A(\read<7> ), .Y(n24) );
  INVX1 U3 ( .A(\read<10> ), .Y(n18) );
  INVX1 U4 ( .A(\read<11> ), .Y(n16) );
  INVX1 U5 ( .A(\read<12> ), .Y(n14) );
  INVX1 U6 ( .A(\read<13> ), .Y(n12) );
  INVX1 U7 ( .A(\read<14> ), .Y(n10) );
  INVX1 U8 ( .A(\read<15> ), .Y(n8) );
  INVX1 U9 ( .A(\read<0> ), .Y(n38) );
  INVX1 U10 ( .A(\read<1> ), .Y(n36) );
  INVX1 U11 ( .A(\read<3> ), .Y(n32) );
  INVX1 U12 ( .A(\read<4> ), .Y(n30) );
  INVX1 U13 ( .A(\read<8> ), .Y(n22) );
  INVX1 U14 ( .A(\read<9> ), .Y(n20) );
  INVX1 U15 ( .A(\read<5> ), .Y(n28) );
  MUX2X1 U16 ( .B(n23), .A(n24), .S(n1), .Y(n46) );
  MUX2X1 U17 ( .B(n7), .A(n8), .S(n4), .Y(n54) );
  INVX1 U18 ( .A(\read<2> ), .Y(n34) );
  INVX1 U19 ( .A(\write<2> ), .Y(n33) );
  INVX1 U20 ( .A(\write<1> ), .Y(n35) );
  INVX1 U21 ( .A(\write<4> ), .Y(n29) );
  BUFX2 U22 ( .A(wr_en), .Y(n6) );
  BUFX2 U23 ( .A(wr_en), .Y(n5) );
  INVX1 U24 ( .A(\write<8> ), .Y(n21) );
  INVX1 U25 ( .A(n6), .Y(n1) );
  MUX2X1 U26 ( .B(n25), .A(n26), .S(n1), .Y(n45) );
  MUX2X1 U27 ( .B(n13), .A(n14), .S(n1), .Y(n51) );
  INVX1 U28 ( .A(\write<5> ), .Y(n27) );
  INVX1 U29 ( .A(\write<3> ), .Y(n31) );
  INVX1 U30 ( .A(\write<0> ), .Y(n37) );
  INVX1 U31 ( .A(\write<12> ), .Y(n13) );
  INVX1 U32 ( .A(\write<6> ), .Y(n25) );
  INVX1 U33 ( .A(\write<9> ), .Y(n19) );
  INVX1 U34 ( .A(n5), .Y(n3) );
  INVX1 U35 ( .A(n5), .Y(n2) );
  INVX1 U36 ( .A(n5), .Y(n4) );
  MUX2X1 U37 ( .B(n11), .A(n12), .S(n2), .Y(n52) );
  INVX1 U38 ( .A(\write<10> ), .Y(n17) );
  INVX1 U39 ( .A(\write<13> ), .Y(n11) );
  INVX1 U40 ( .A(\write<7> ), .Y(n23) );
  MUX2X1 U41 ( .B(n9), .A(n10), .S(n3), .Y(n53) );
  INVX1 U42 ( .A(\write<14> ), .Y(n9) );
  MUX2X1 U43 ( .B(n15), .A(n16), .S(n4), .Y(n50) );
  INVX1 U44 ( .A(\write<15> ), .Y(n7) );
  INVX1 U45 ( .A(\write<11> ), .Y(n15) );
  MUX2X1 U46 ( .B(n18), .A(n17), .S(n6), .Y(n49) );
  MUX2X1 U47 ( .B(n20), .A(n19), .S(n5), .Y(n48) );
  MUX2X1 U48 ( .B(n22), .A(n21), .S(n5), .Y(n47) );
  MUX2X1 U49 ( .B(n28), .A(n27), .S(n6), .Y(n44) );
  MUX2X1 U50 ( .B(n30), .A(n29), .S(n6), .Y(n43) );
  MUX2X1 U51 ( .B(n32), .A(n31), .S(n5), .Y(n42) );
  MUX2X1 U52 ( .B(n34), .A(n33), .S(n5), .Y(n41) );
  MUX2X1 U53 ( .B(n36), .A(n35), .S(n5), .Y(n40) );
  MUX2X1 U54 ( .B(n38), .A(n37), .S(n6), .Y(n39) );
endmodule


module CLA16_5 ( .A({\A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , 
        \A<9> , \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , 
        \A<0> }), .B({\B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , 
        \B<9> , \B<8> , \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , 
        \B<0> }), Cin, Cout, .S({\S<15> , \S<14> , \S<13> , \S<12> , \S<11> , 
        \S<10> , \S<9> , \S<8> , \S<7> , \S<6> , \S<5> , \S<4> , \S<3> , 
        \S<2> , \S<1> , \S<0> }) );
  input \A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> , \A<8> ,
         \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , \A<0> ,
         \B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , \B<9> , \B<8> ,
         \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output Cout, \S<15> , \S<14> , \S<13> , \S<12> , \S<11> , \S<10> , \S<9> ,
         \S<8> , \S<7> , \S<6> , \S<5> , \S<4> , \S<3> , \S<2> , \S<1> ,
         \S<0> ;
  wire   p30, g30, p74, g74, p118, g118, p1512, g1512, n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22;

  CLA4_23 A3_0 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), .Cin(Cin), .Cout(), .P(p30), .G(g30), .S({\S<3> , 
        \S<2> , \S<1> , \S<0> }) );
  CLA4_22 A7_4 ( .A({\A<7> , \A<6> , \A<5> , \A<4> }), .B({\B<7> , \B<6> , 
        \B<5> , \B<4> }), .Cin(n3), .Cout(), .P(p74), .G(g74), .S({\S<7> , 
        \S<6> , \S<5> , \S<4> }) );
  CLA4_21 A11_8 ( .A({\A<11> , \A<10> , \A<9> , \A<8> }), .B({\B<11> , \B<10> , 
        \B<9> , \B<8> }), .Cin(n6), .Cout(), .P(p118), .G(g118), .S({\S<11> , 
        \S<10> , \S<9> , \S<8> }) );
  CLA4_20 A15_12 ( .A({\A<15> , \A<14> , \A<13> , \A<12> }), .B({\B<15> , 
        \B<14> , \B<13> , \B<12> }), .Cin(n13), .Cout(), .P(p1512), .G(g1512), 
        .S({\S<15> , \S<14> , \S<13> , \S<12> }) );
  INVX1 U1 ( .A(g1512), .Y(n21) );
  INVX1 U2 ( .A(p1512), .Y(n22) );
  INVX1 U3 ( .A(g118), .Y(n20) );
  AND2X2 U4 ( .A(p118), .B(n6), .Y(n11) );
  INVX1 U5 ( .A(g30), .Y(n1) );
  INVX2 U6 ( .A(n2), .Y(n3) );
  AND2X2 U7 ( .A(n1), .B(n10), .Y(n2) );
  AND2X2 U8 ( .A(n18), .B(n17), .Y(n4) );
  INVX1 U9 ( .A(n4), .Y(n5) );
  AND2X2 U10 ( .A(n15), .B(n5), .Y(n6) );
  OR2X1 U11 ( .A(n16), .B(p74), .Y(n15) );
  INVX1 U12 ( .A(n10), .Y(n7) );
  INVX1 U13 ( .A(n7), .Y(n8) );
  AND2X1 U14 ( .A(Cin), .B(p30), .Y(n9) );
  INVX1 U15 ( .A(n9), .Y(n10) );
  INVX1 U16 ( .A(n11), .Y(n12) );
  INVX1 U17 ( .A(n14), .Y(n13) );
  AND2X2 U18 ( .A(n20), .B(n12), .Y(n14) );
  INVX1 U19 ( .A(g74), .Y(n19) );
  INVX1 U20 ( .A(g30), .Y(n18) );
  INVX1 U21 ( .A(n19), .Y(n16) );
  AND2X2 U22 ( .A(n8), .B(n19), .Y(n17) );
  OAI21X1 U23 ( .A(n14), .B(n22), .C(n21), .Y(Cout) );
endmodule


module CLA16_4 ( .A({\A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , 
        \A<9> , \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , 
        \A<0> }), .B({\B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , 
        \B<9> , \B<8> , \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , 
        \B<0> }), Cin, Cout, .S({\S<15> , \S<14> , \S<13> , \S<12> , \S<11> , 
        \S<10> , \S<9> , \S<8> , \S<7> , \S<6> , \S<5> , \S<4> , \S<3> , 
        \S<2> , \S<1> , \S<0> }) );
  input \A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> , \A<8> ,
         \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , \A<0> ,
         \B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , \B<9> , \B<8> ,
         \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output Cout, \S<15> , \S<14> , \S<13> , \S<12> , \S<11> , \S<10> , \S<9> ,
         \S<8> , \S<7> , \S<6> , \S<5> , \S<4> , \S<3> , \S<2> , \S<1> ,
         \S<0> ;
  wire   p30, g30, p74, g74, p118, g118, p1512, g1512, n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n14, n15;

  CLA4_19 A3_0 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), .Cin(Cin), .Cout(), .P(p30), .G(g30), .S({\S<3> , 
        \S<2> , \S<1> , \S<0> }) );
  CLA4_18 A7_4 ( .A({\A<7> , \A<6> , \A<5> , \A<4> }), .B({\B<7> , \B<6> , 
        \B<5> , \B<4> }), .Cin(n15), .Cout(), .P(p74), .G(g74), .S({\S<7> , 
        \S<6> , \S<5> , \S<4> }) );
  CLA4_17 A11_8 ( .A({\A<11> , \A<10> , \A<9> , \A<8> }), .B({\B<11> , \B<10> , 
        \B<9> , \B<8> }), .Cin(n14), .Cout(), .P(p118), .G(g118), .S({\S<11> , 
        \S<10> , \S<9> , \S<8> }) );
  CLA4_16 A15_12 ( .A({\A<15> , \A<14> , \A<13> , \A<12> }), .B({\B<15> , 
        \B<14> , \B<13> , \B<12> }), .Cin(n5), .Cout(), .P(p1512), .G(g1512), 
        .S({\S<15> , \S<14> , \S<13> , \S<12> }) );
  INVX1 U1 ( .A(g118), .Y(n9) );
  INVX1 U2 ( .A(g1512), .Y(n10) );
  INVX1 U3 ( .A(p1512), .Y(n11) );
  INVX1 U4 ( .A(n5), .Y(n12) );
  INVX1 U5 ( .A(n4), .Y(n14) );
  INVX2 U6 ( .A(n6), .Y(n5) );
  INVX2 U7 ( .A(n1), .Y(n15) );
  BUFX2 U8 ( .A(n8), .Y(n1) );
  AND2X2 U9 ( .A(p118), .B(n14), .Y(n2) );
  INVX1 U10 ( .A(n2), .Y(n3) );
  BUFX2 U11 ( .A(n7), .Y(n4) );
  AND2X2 U12 ( .A(n9), .B(n3), .Y(n6) );
  AOI21X1 U13 ( .A(n15), .B(p74), .C(g74), .Y(n7) );
  AOI21X1 U14 ( .A(Cin), .B(p30), .C(g30), .Y(n8) );
  OAI21X1 U15 ( .A(n12), .B(n11), .C(n10), .Y(Cout) );
endmodule


module CLA16_3 ( .A({\A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , 
        \A<9> , \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , 
        \A<0> }), .B({\B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , 
        \B<9> , \B<8> , \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , 
        \B<0> }), Cin, Cout, .S({\S<15> , \S<14> , \S<13> , \S<12> , \S<11> , 
        \S<10> , \S<9> , \S<8> , \S<7> , \S<6> , \S<5> , \S<4> , \S<3> , 
        \S<2> , \S<1> , \S<0> }) );
  input \A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> , \A<8> ,
         \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , \A<0> ,
         \B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , \B<9> , \B<8> ,
         \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output Cout, \S<15> , \S<14> , \S<13> , \S<12> , \S<11> , \S<10> , \S<9> ,
         \S<8> , \S<7> , \S<6> , \S<5> , \S<4> , \S<3> , \S<2> , \S<1> ,
         \S<0> ;
  wire   p30, g30, p74, g74, p118, g118, p1512, g1512, n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n19;

  CLA4_15 A3_0 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), .Cin(Cin), .Cout(), .P(p30), .G(g30), .S({\S<3> , 
        \S<2> , \S<1> , \S<0> }) );
  CLA4_14 A7_4 ( .A({\A<7> , \A<6> , \A<5> , \A<4> }), .B({\B<7> , \B<6> , 
        \B<5> , \B<4> }), .Cin(n7), .Cout(), .P(p74), .G(g74), .S({\S<7> , 
        \S<6> , \S<5> , \S<4> }) );
  CLA4_13 A11_8 ( .A({\A<11> , \A<10> , \A<9> , \A<8> }), .B({\B<11> , \B<10> , 
        \B<9> , \B<8> }), .Cin(n3), .Cout(), .P(p118), .G(g118), .S({\S<11> , 
        \S<10> , \S<9> , \S<8> }) );
  CLA4_12 A15_12 ( .A({\A<15> , \A<14> , \A<13> , \A<12> }), .B({\B<15> , 
        \B<14> , \B<13> , \B<12> }), .Cin(n1), .Cout(), .P(p1512), .G(g1512), 
        .S({\S<15> , \S<14> , \S<13> , \S<12> }) );
  INVX1 U1 ( .A(p1512), .Y(n17) );
  INVX1 U2 ( .A(n10), .Y(n1) );
  INVX1 U3 ( .A(n5), .Y(n12) );
  AND2X2 U4 ( .A(n14), .B(n13), .Y(n10) );
  AND2X2 U5 ( .A(n15), .B(n8), .Y(n2) );
  INVX1 U6 ( .A(n2), .Y(n3) );
  AND2X2 U7 ( .A(p74), .B(n19), .Y(n4) );
  INVX1 U8 ( .A(n4), .Y(n5) );
  INVX1 U9 ( .A(n19), .Y(n6) );
  INVX1 U10 ( .A(n6), .Y(n7) );
  INVX1 U11 ( .A(n11), .Y(n19) );
  INVX1 U12 ( .A(g1512), .Y(n16) );
  INVX1 U13 ( .A(g74), .Y(n15) );
  INVX1 U14 ( .A(n4), .Y(n8) );
  INVX1 U15 ( .A(n1), .Y(n9) );
  INVX1 U16 ( .A(g118), .Y(n14) );
  AOI21X1 U17 ( .A(Cin), .B(p30), .C(g30), .Y(n11) );
  OAI21X1 U18 ( .A(n12), .B(g74), .C(p118), .Y(n13) );
  OAI21X1 U19 ( .A(n9), .B(n17), .C(n16), .Y(Cout) );
endmodule


module CLA16_2 ( .A({\A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , 
        \A<9> , \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , 
        \A<0> }), .B({\B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , 
        \B<9> , \B<8> , \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , 
        \B<0> }), Cin, Cout, .S({\S<15> , \S<14> , \S<13> , \S<12> , \S<11> , 
        \S<10> , \S<9> , \S<8> , \S<7> , \S<6> , \S<5> , \S<4> , \S<3> , 
        \S<2> , \S<1> , \S<0> }) );
  input \A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> , \A<8> ,
         \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , \A<0> ,
         \B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , \B<9> , \B<8> ,
         \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output Cout, \S<15> , \S<14> , \S<13> , \S<12> , \S<11> , \S<10> , \S<9> ,
         \S<8> , \S<7> , \S<6> , \S<5> , \S<4> , \S<3> , \S<2> , \S<1> ,
         \S<0> ;
  wire   p30, g30, p74, g74, p118, g118, p1512, g1512, n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n16, n17;

  CLA4_11 A3_0 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), .Cin(Cin), .Cout(), .P(p30), .G(g30), .S({\S<3> , 
        \S<2> , \S<1> , \S<0> }) );
  CLA4_10 A7_4 ( .A({\A<7> , \A<6> , \A<5> , \A<4> }), .B({\B<7> , \B<6> , 
        \B<5> , \B<4> }), .Cin(n17), .Cout(), .P(p74), .G(g74), .S({\S<7> , 
        \S<6> , \S<5> , \S<4> }) );
  CLA4_9 A11_8 ( .A({\A<11> , \A<10> , \A<9> , \A<8> }), .B({\B<11> , \B<10> , 
        \B<9> , \B<8> }), .Cin(n3), .Cout(), .P(p118), .G(g118), .S({\S<11> , 
        \S<10> , \S<9> , \S<8> }) );
  CLA4_8 A15_12 ( .A({\A<15> , \A<14> , \A<13> , \A<12> }), .B({\B<15> , 
        \B<14> , \B<13> , \B<12> }), .Cin(n16), .Cout(), .P(p1512), .G(g1512), 
        .S({\S<15> , \S<14> , \S<13> , \S<12> }) );
  INVX1 U1 ( .A(g1512), .Y(n13) );
  INVX1 U2 ( .A(n12), .Y(n1) );
  INVX4 U3 ( .A(n7), .Y(n16) );
  AND2X2 U4 ( .A(n12), .B(n4), .Y(n2) );
  INVX1 U5 ( .A(n2), .Y(n3) );
  INVX1 U6 ( .A(n6), .Y(n4) );
  AND2X2 U7 ( .A(p74), .B(n17), .Y(n6) );
  BUFX2 U8 ( .A(n8), .Y(n5) );
  INVX1 U9 ( .A(p1512), .Y(n14) );
  INVX1 U10 ( .A(g74), .Y(n12) );
  INVX1 U11 ( .A(n4), .Y(n9) );
  AND2X2 U12 ( .A(n11), .B(n10), .Y(n7) );
  INVX1 U13 ( .A(g118), .Y(n11) );
  AOI21X1 U14 ( .A(Cin), .B(p30), .C(g30), .Y(n8) );
  INVX2 U15 ( .A(n5), .Y(n17) );
  OAI21X1 U16 ( .A(n1), .B(n9), .C(p118), .Y(n10) );
  OAI21X1 U17 ( .A(n7), .B(n14), .C(n13), .Y(Cout) );
endmodule


module CLA16_1 ( .A({\A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , 
        \A<9> , \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , 
        \A<0> }), .B({\B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , 
        \B<9> , \B<8> , \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , 
        \B<0> }), Cin, Cout, .S({\S<15> , \S<14> , \S<13> , \S<12> , \S<11> , 
        \S<10> , \S<9> , \S<8> , \S<7> , \S<6> , \S<5> , \S<4> , \S<3> , 
        \S<2> , \S<1> , \S<0> }) );
  input \A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> , \A<8> ,
         \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , \A<0> ,
         \B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , \B<9> , \B<8> ,
         \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output Cout, \S<15> , \S<14> , \S<13> , \S<12> , \S<11> , \S<10> , \S<9> ,
         \S<8> , \S<7> , \S<6> , \S<5> , \S<4> , \S<3> , \S<2> , \S<1> ,
         \S<0> ;
  wire   p30, g30, p74, g74, p118, g118, p1512, g1512, n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14;

  CLA4_7 A3_0 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), .Cin(Cin), .Cout(), .P(p30), .G(g30), .S({\S<3> , 
        \S<2> , \S<1> , \S<0> }) );
  CLA4_6 A7_4 ( .A({\A<7> , \A<6> , \A<5> , \A<4> }), .B({\B<7> , \B<6> , 
        \B<5> , \B<4> }), .Cin(n3), .Cout(), .P(p74), .G(g74), .S({\S<7> , 
        \S<6> , \S<5> , \S<4> }) );
  CLA4_5 A11_8 ( .A({\A<11> , \A<10> , \A<9> , \A<8> }), .B({\B<11> , \B<10> , 
        \B<9> , \B<8> }), .Cin(n14), .Cout(), .P(p118), .G(g118), .S({\S<11> , 
        \S<10> , \S<9> , \S<8> }) );
  CLA4_4 A15_12 ( .A({\A<15> , \A<14> , \A<13> , \A<12> }), .B({\B<15> , 
        \B<14> , \B<13> , \B<12> }), .Cin(n1), .Cout(), .P(p1512), .G(g1512), 
        .S({\S<15> , \S<14> , \S<13> , \S<12> }) );
  INVX1 U1 ( .A(g1512), .Y(n12) );
  INVX1 U2 ( .A(p1512), .Y(n13) );
  INVX1 U3 ( .A(p74), .Y(n11) );
  INVX1 U4 ( .A(g74), .Y(n10) );
  OR2X2 U5 ( .A(n7), .B(g118), .Y(n1) );
  AND2X2 U6 ( .A(n5), .B(n8), .Y(n2) );
  INVX1 U7 ( .A(n2), .Y(n3) );
  AND2X2 U8 ( .A(Cin), .B(p30), .Y(n4) );
  INVX1 U9 ( .A(n4), .Y(n5) );
  INVX1 U10 ( .A(n1), .Y(n6) );
  AND2X2 U11 ( .A(n9), .B(p118), .Y(n7) );
  INVX1 U12 ( .A(g30), .Y(n8) );
  OAI21X1 U13 ( .A(n11), .B(n2), .C(n10), .Y(n9) );
  OAI21X1 U14 ( .A(n2), .B(n11), .C(n10), .Y(n14) );
  OAI21X1 U15 ( .A(n6), .B(n13), .C(n12), .Y(Cout) );
endmodule


module dff_647 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_646 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_645 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_644 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_643 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_642 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X1 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_641 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_640 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_639 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_638 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_637 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_636 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_635 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_634 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_633 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_632 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_631 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_630 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_629 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_628 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_627 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_626 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_625 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_624 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_623 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_622 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_621 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_620 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_619 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_618 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_617 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_616 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_615 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_614 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_613 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_612 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_611 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_610 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_609 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_608 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_607 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_606 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_605 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_604 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_603 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_602 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_601 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_600 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_599 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_598 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module rf ( .read1data({\read1data<15> , \read1data<14> , \read1data<13> , 
        \read1data<12> , \read1data<11> , \read1data<10> , \read1data<9> , 
        \read1data<8> , \read1data<7> , \read1data<6> , \read1data<5> , 
        \read1data<4> , \read1data<3> , \read1data<2> , \read1data<1> , 
        \read1data<0> }), .read2data({\read2data<15> , \read2data<14> , 
        \read2data<13> , \read2data<12> , \read2data<11> , \read2data<10> , 
        \read2data<9> , \read2data<8> , \read2data<7> , \read2data<6> , 
        \read2data<5> , \read2data<4> , \read2data<3> , \read2data<2> , 
        \read2data<1> , \read2data<0> }), err, clk, rst, .read1regsel({
        \read1regsel<2> , \read1regsel<1> , \read1regsel<0> }), .read2regsel({
        \read2regsel<2> , \read2regsel<1> , \read2regsel<0> }), .writeregsel({
        \writeregsel<2> , \writeregsel<1> , \writeregsel<0> }), .writedata({
        \writedata<15> , \writedata<14> , \writedata<13> , \writedata<12> , 
        \writedata<11> , \writedata<10> , \writedata<9> , \writedata<8> , 
        \writedata<7> , \writedata<6> , \writedata<5> , \writedata<4> , 
        \writedata<3> , \writedata<2> , \writedata<1> , \writedata<0> }), 
        write );
  input clk, rst, \read1regsel<2> , \read1regsel<1> , \read1regsel<0> ,
         \read2regsel<2> , \read2regsel<1> , \read2regsel<0> ,
         \writeregsel<2> , \writeregsel<1> , \writeregsel<0> , \writedata<15> ,
         \writedata<14> , \writedata<13> , \writedata<12> , \writedata<11> ,
         \writedata<10> , \writedata<9> , \writedata<8> , \writedata<7> ,
         \writedata<6> , \writedata<5> , \writedata<4> , \writedata<3> ,
         \writedata<2> , \writedata<1> , \writedata<0> , write;
  output \read1data<15> , \read1data<14> , \read1data<13> , \read1data<12> ,
         \read1data<11> , \read1data<10> , \read1data<9> , \read1data<8> ,
         \read1data<7> , \read1data<6> , \read1data<5> , \read1data<4> ,
         \read1data<3> , \read1data<2> , \read1data<1> , \read1data<0> ,
         \read2data<15> , \read2data<14> , \read2data<13> , \read2data<12> ,
         \read2data<11> , \read2data<10> , \read2data<9> , \read2data<8> ,
         \read2data<7> , \read2data<6> , \read2data<5> , \read2data<4> ,
         \read2data<3> , \read2data<2> , \read2data<1> , \read2data<0> , err;
  wire   n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         \writedecode<7> , \writedecode<6> , \writedecode<5> ,
         \writedecode<4> , \writedecode<3> , \writedecode<2> ,
         \writedecode<1> , \writedecode<0> , \readoutR0<15> , \readoutR0<14> ,
         \readoutR0<13> , \readoutR0<12> , \readoutR0<11> , \readoutR0<10> ,
         \readoutR0<9> , \readoutR0<8> , \readoutR0<7> , \readoutR0<6> ,
         \readoutR0<5> , \readoutR0<4> , \readoutR0<3> , \readoutR0<2> ,
         \readoutR0<1> , \readoutR0<0> , \readoutR1<15> , \readoutR1<14> ,
         \readoutR1<13> , \readoutR1<12> , \readoutR1<11> , \readoutR1<10> ,
         \readoutR1<9> , \readoutR1<8> , \readoutR1<7> , \readoutR1<6> ,
         \readoutR1<5> , \readoutR1<4> , \readoutR1<3> , \readoutR1<2> ,
         \readoutR1<1> , \readoutR1<0> , \readoutR2<15> , \readoutR2<14> ,
         \readoutR2<13> , \readoutR2<12> , \readoutR2<11> , \readoutR2<10> ,
         \readoutR2<9> , \readoutR2<8> , \readoutR2<7> , \readoutR2<6> ,
         \readoutR2<5> , \readoutR2<4> , \readoutR2<3> , \readoutR2<2> ,
         \readoutR2<1> , \readoutR2<0> , \readoutR3<15> , \readoutR3<14> ,
         \readoutR3<13> , \readoutR3<12> , \readoutR3<11> , \readoutR3<10> ,
         \readoutR3<9> , \readoutR3<8> , \readoutR3<7> , \readoutR3<6> ,
         \readoutR3<5> , \readoutR3<4> , \readoutR3<3> , \readoutR3<2> ,
         \readoutR3<1> , \readoutR3<0> , \readoutR4<15> , \readoutR4<14> ,
         \readoutR4<13> , \readoutR4<12> , \readoutR4<11> , \readoutR4<10> ,
         \readoutR4<9> , \readoutR4<8> , \readoutR4<7> , \readoutR4<6> ,
         \readoutR4<5> , \readoutR4<4> , \readoutR4<3> , \readoutR4<2> ,
         \readoutR4<1> , \readoutR4<0> , \readoutR5<15> , \readoutR5<14> ,
         \readoutR5<13> , \readoutR5<12> , \readoutR5<11> , \readoutR5<10> ,
         \readoutR5<9> , \readoutR5<8> , \readoutR5<7> , \readoutR5<6> ,
         \readoutR5<5> , \readoutR5<4> , \readoutR5<3> , \readoutR5<2> ,
         \readoutR5<1> , \readoutR5<0> , \readoutR6<15> , \readoutR6<14> ,
         \readoutR6<13> , \readoutR6<12> , \readoutR6<11> , \readoutR6<10> ,
         \readoutR6<9> , \readoutR6<8> , \readoutR6<7> , \readoutR6<6> ,
         \readoutR6<5> , \readoutR6<4> , \readoutR6<3> , \readoutR6<2> ,
         \readoutR6<1> , \readoutR6<0> , \readoutR7<15> , \readoutR7<14> ,
         \readoutR7<13> , \readoutR7<12> , \readoutR7<11> , \readoutR7<10> ,
         \readoutR7<9> , \readoutR7<8> , \readoutR7<7> , \readoutR7<6> ,
         \readoutR7<5> , \readoutR7<4> , \readoutR7<3> , \readoutR7<2> ,
         \readoutR7<1> , \readoutR7<0> , n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n1, n17, n18,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n306, n308, n310, n312, n314, n316, n318, n320, n322, n324, n326,
         n328, n330, n332, n334, n336, n338, n340, n342, n344, n346, n348,
         n350, n352, n354, n356, n358, n360, n362, n364, n366, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451;
  assign err = 1'b0;

  reg16_7 r0 ( .read({\readoutR0<15> , \readoutR0<14> , \readoutR0<13> , 
        \readoutR0<12> , \readoutR0<11> , \readoutR0<10> , \readoutR0<9> , 
        \readoutR0<8> , \readoutR0<7> , \readoutR0<6> , \readoutR0<5> , 
        \readoutR0<4> , \readoutR0<3> , \readoutR0<2> , \readoutR0<1> , 
        \readoutR0<0> }), .write({\writedata<15> , \writedata<14> , 
        \writedata<13> , \writedata<12> , \writedata<11> , \writedata<10> , 
        \writedata<9> , \writedata<8> , \writedata<7> , \writedata<6> , 
        \writedata<5> , \writedata<4> , \writedata<3> , \writedata<2> , 
        \writedata<1> , \writedata<0> }), .wr_en(\writedecode<0> ), .rst(rst), 
        .clk(clk) );
  reg16_6 r1 ( .read({\readoutR1<15> , \readoutR1<14> , \readoutR1<13> , 
        \readoutR1<12> , \readoutR1<11> , \readoutR1<10> , \readoutR1<9> , 
        \readoutR1<8> , \readoutR1<7> , \readoutR1<6> , \readoutR1<5> , 
        \readoutR1<4> , \readoutR1<3> , \readoutR1<2> , \readoutR1<1> , 
        \readoutR1<0> }), .write({\writedata<15> , \writedata<14> , 
        \writedata<13> , \writedata<12> , \writedata<11> , \writedata<10> , 
        \writedata<9> , \writedata<8> , \writedata<7> , \writedata<6> , 
        \writedata<5> , \writedata<4> , \writedata<3> , \writedata<2> , 
        \writedata<1> , \writedata<0> }), .wr_en(\writedecode<1> ), .rst(rst), 
        .clk(clk) );
  reg16_5 r2 ( .read({\readoutR2<15> , \readoutR2<14> , \readoutR2<13> , 
        \readoutR2<12> , \readoutR2<11> , \readoutR2<10> , \readoutR2<9> , 
        \readoutR2<8> , \readoutR2<7> , \readoutR2<6> , \readoutR2<5> , 
        \readoutR2<4> , \readoutR2<3> , \readoutR2<2> , \readoutR2<1> , 
        \readoutR2<0> }), .write({\writedata<15> , \writedata<14> , 
        \writedata<13> , \writedata<12> , \writedata<11> , \writedata<10> , 
        \writedata<9> , \writedata<8> , \writedata<7> , \writedata<6> , 
        \writedata<5> , \writedata<4> , \writedata<3> , \writedata<2> , 
        \writedata<1> , \writedata<0> }), .wr_en(\writedecode<2> ), .rst(rst), 
        .clk(clk) );
  reg16_4 r3 ( .read({\readoutR3<15> , \readoutR3<14> , \readoutR3<13> , 
        \readoutR3<12> , \readoutR3<11> , \readoutR3<10> , \readoutR3<9> , 
        \readoutR3<8> , \readoutR3<7> , \readoutR3<6> , \readoutR3<5> , 
        \readoutR3<4> , \readoutR3<3> , \readoutR3<2> , \readoutR3<1> , 
        \readoutR3<0> }), .write({\writedata<15> , \writedata<14> , 
        \writedata<13> , \writedata<12> , \writedata<11> , \writedata<10> , 
        \writedata<9> , \writedata<8> , \writedata<7> , \writedata<6> , 
        \writedata<5> , \writedata<4> , \writedata<3> , \writedata<2> , 
        \writedata<1> , \writedata<0> }), .wr_en(\writedecode<3> ), .rst(rst), 
        .clk(clk) );
  reg16_3 r4 ( .read({\readoutR4<15> , \readoutR4<14> , \readoutR4<13> , 
        \readoutR4<12> , \readoutR4<11> , \readoutR4<10> , \readoutR4<9> , 
        \readoutR4<8> , \readoutR4<7> , \readoutR4<6> , \readoutR4<5> , 
        \readoutR4<4> , \readoutR4<3> , \readoutR4<2> , \readoutR4<1> , 
        \readoutR4<0> }), .write({\writedata<15> , \writedata<14> , 
        \writedata<13> , \writedata<12> , \writedata<11> , \writedata<10> , 
        \writedata<9> , \writedata<8> , \writedata<7> , \writedata<6> , 
        \writedata<5> , \writedata<4> , \writedata<3> , \writedata<2> , 
        \writedata<1> , \writedata<0> }), .wr_en(\writedecode<4> ), .rst(rst), 
        .clk(clk) );
  reg16_2 r5 ( .read({\readoutR5<15> , \readoutR5<14> , \readoutR5<13> , 
        \readoutR5<12> , \readoutR5<11> , \readoutR5<10> , \readoutR5<9> , 
        \readoutR5<8> , \readoutR5<7> , \readoutR5<6> , \readoutR5<5> , 
        \readoutR5<4> , \readoutR5<3> , \readoutR5<2> , \readoutR5<1> , 
        \readoutR5<0> }), .write({\writedata<15> , \writedata<14> , 
        \writedata<13> , \writedata<12> , \writedata<11> , \writedata<10> , 
        \writedata<9> , \writedata<8> , \writedata<7> , \writedata<6> , 
        \writedata<5> , \writedata<4> , \writedata<3> , \writedata<2> , 
        \writedata<1> , \writedata<0> }), .wr_en(\writedecode<5> ), .rst(rst), 
        .clk(clk) );
  reg16_1 r6 ( .read({\readoutR6<15> , \readoutR6<14> , \readoutR6<13> , 
        \readoutR6<12> , \readoutR6<11> , \readoutR6<10> , \readoutR6<9> , 
        \readoutR6<8> , \readoutR6<7> , \readoutR6<6> , \readoutR6<5> , 
        \readoutR6<4> , \readoutR6<3> , \readoutR6<2> , \readoutR6<1> , 
        \readoutR6<0> }), .write({\writedata<15> , \writedata<14> , 
        \writedata<13> , \writedata<12> , \writedata<11> , \writedata<10> , 
        \writedata<9> , \writedata<8> , \writedata<7> , \writedata<6> , 
        \writedata<5> , \writedata<4> , \writedata<3> , \writedata<2> , 
        \writedata<1> , \writedata<0> }), .wr_en(\writedecode<6> ), .rst(rst), 
        .clk(clk) );
  reg16_0 r7 ( .read({\readoutR7<15> , \readoutR7<14> , \readoutR7<13> , 
        \readoutR7<12> , \readoutR7<11> , \readoutR7<10> , \readoutR7<9> , 
        \readoutR7<8> , \readoutR7<7> , \readoutR7<6> , \readoutR7<5> , 
        \readoutR7<4> , \readoutR7<3> , \readoutR7<2> , \readoutR7<1> , 
        \readoutR7<0> }), .write({\writedata<15> , \writedata<14> , 
        \writedata<13> , \writedata<12> , \writedata<11> , \writedata<10> , 
        \writedata<9> , \writedata<8> , \writedata<7> , \writedata<6> , 
        \writedata<5> , \writedata<4> , \writedata<3> , \writedata<2> , 
        \writedata<1> , \writedata<0> }), .wr_en(\writedecode<7> ), .rst(rst), 
        .clk(clk) );
  AND2X2 U2 ( .A(n255), .B(n271), .Y(n21) );
  AND2X2 U3 ( .A(n253), .B(n270), .Y(n30) );
  AND2X2 U4 ( .A(n251), .B(n269), .Y(n35) );
  AND2X2 U5 ( .A(n249), .B(n268), .Y(n40) );
  AND2X2 U6 ( .A(n247), .B(n267), .Y(n45) );
  AND2X2 U7 ( .A(n245), .B(n266), .Y(n50) );
  AND2X2 U8 ( .A(n243), .B(n265), .Y(n55) );
  AND2X2 U9 ( .A(n241), .B(n264), .Y(n60) );
  AND2X2 U10 ( .A(n239), .B(n263), .Y(n65) );
  AND2X2 U11 ( .A(n237), .B(n262), .Y(n70) );
  AND2X2 U12 ( .A(n235), .B(n261), .Y(n75) );
  AND2X2 U13 ( .A(n233), .B(n260), .Y(n80) );
  AND2X2 U14 ( .A(n231), .B(n259), .Y(n85) );
  AND2X2 U15 ( .A(n229), .B(n258), .Y(n90) );
  AND2X2 U16 ( .A(n227), .B(n257), .Y(n95) );
  AND2X2 U17 ( .A(n225), .B(n256), .Y(n100) );
  INVX2 U38 ( .A(\read1regsel<1> ), .Y(n6) );
  INVX2 U39 ( .A(\read1regsel<0> ), .Y(n7) );
  INVX2 U45 ( .A(\read2regsel<0> ), .Y(n13) );
  NOR3X1 U49 ( .A(n14), .B(n443), .C(n15), .Y(\writedecode<7> ) );
  NOR3X1 U50 ( .A(n441), .B(n15), .C(n14), .Y(\writedecode<6> ) );
  NOR3X1 U51 ( .A(n14), .B(\writeregsel<1> ), .C(n443), .Y(\writedecode<5> )
         );
  NOR3X1 U52 ( .A(n441), .B(\writeregsel<1> ), .C(n14), .Y(\writedecode<4> )
         );
  NOR3X1 U53 ( .A(n15), .B(\writeregsel<2> ), .C(n443), .Y(\writedecode<3> )
         );
  NOR3X1 U54 ( .A(n441), .B(\writeregsel<2> ), .C(n15), .Y(\writedecode<2> )
         );
  NOR3X1 U55 ( .A(n443), .B(\writeregsel<2> ), .C(\writeregsel<1> ), .Y(
        \writedecode<1> ) );
  NOR3X1 U57 ( .A(n441), .B(\writeregsel<2> ), .C(\writeregsel<1> ), .Y(
        \writedecode<0> ) );
  NAND3X1 U59 ( .A(n399), .B(n431), .C(n21), .Y(n474) );
  AOI22X1 U60 ( .A(\readoutR7<9> ), .B(n9), .C(\readoutR6<9> ), .D(n8), .Y(n23) );
  AOI22X1 U61 ( .A(\readoutR5<9> ), .B(n11), .C(\readoutR4<9> ), .D(n10), .Y(
        n22) );
  AOI22X1 U62 ( .A(\readoutR3<9> ), .B(n450), .C(\readoutR2<9> ), .D(n451), 
        .Y(n20) );
  AOI22X1 U63 ( .A(\readoutR1<9> ), .B(n448), .C(\readoutR0<9> ), .D(n449), 
        .Y(n19) );
  NAND3X1 U64 ( .A(n398), .B(n430), .C(n30), .Y(n475) );
  AOI22X1 U65 ( .A(\readoutR7<8> ), .B(n9), .C(\readoutR6<8> ), .D(n8), .Y(n32) );
  AOI22X1 U66 ( .A(\readoutR5<8> ), .B(n11), .C(\readoutR4<8> ), .D(n10), .Y(
        n31) );
  AOI22X1 U67 ( .A(\readoutR3<8> ), .B(n450), .C(\readoutR2<8> ), .D(n451), 
        .Y(n29) );
  AOI22X1 U68 ( .A(\readoutR1<8> ), .B(n448), .C(\readoutR0<8> ), .D(n449), 
        .Y(n28) );
  NAND3X1 U69 ( .A(n397), .B(n429), .C(n35), .Y(n476) );
  AOI22X1 U70 ( .A(\readoutR7<7> ), .B(n9), .C(\readoutR6<7> ), .D(n8), .Y(n37) );
  AOI22X1 U71 ( .A(\readoutR5<7> ), .B(n11), .C(\readoutR4<7> ), .D(n10), .Y(
        n36) );
  AOI22X1 U72 ( .A(\readoutR3<7> ), .B(n450), .C(\readoutR2<7> ), .D(n451), 
        .Y(n34) );
  AOI22X1 U73 ( .A(\readoutR1<7> ), .B(n448), .C(\readoutR0<7> ), .D(n449), 
        .Y(n33) );
  NAND3X1 U74 ( .A(n396), .B(n428), .C(n40), .Y(n477) );
  AOI22X1 U75 ( .A(\readoutR7<6> ), .B(n9), .C(\readoutR6<6> ), .D(n8), .Y(n42) );
  AOI22X1 U76 ( .A(\readoutR5<6> ), .B(n11), .C(\readoutR4<6> ), .D(n10), .Y(
        n41) );
  AOI22X1 U77 ( .A(\readoutR3<6> ), .B(n450), .C(\readoutR2<6> ), .D(n451), 
        .Y(n39) );
  AOI22X1 U78 ( .A(\readoutR1<6> ), .B(n448), .C(\readoutR0<6> ), .D(n449), 
        .Y(n38) );
  NAND3X1 U79 ( .A(n395), .B(n427), .C(n45), .Y(n478) );
  AOI22X1 U80 ( .A(\readoutR7<5> ), .B(n9), .C(\readoutR6<5> ), .D(n8), .Y(n47) );
  AOI22X1 U81 ( .A(\readoutR5<5> ), .B(n11), .C(\readoutR4<5> ), .D(n10), .Y(
        n46) );
  AOI22X1 U82 ( .A(\readoutR3<5> ), .B(n450), .C(\readoutR2<5> ), .D(n451), 
        .Y(n44) );
  AOI22X1 U83 ( .A(\readoutR1<5> ), .B(n448), .C(\readoutR0<5> ), .D(n449), 
        .Y(n43) );
  NAND3X1 U84 ( .A(n394), .B(n426), .C(n50), .Y(n479) );
  AOI22X1 U85 ( .A(\readoutR7<4> ), .B(n9), .C(\readoutR6<4> ), .D(n8), .Y(n52) );
  AOI22X1 U86 ( .A(\readoutR5<4> ), .B(n11), .C(\readoutR4<4> ), .D(n10), .Y(
        n51) );
  AOI22X1 U87 ( .A(\readoutR3<4> ), .B(n450), .C(\readoutR2<4> ), .D(n451), 
        .Y(n49) );
  AOI22X1 U88 ( .A(\readoutR1<4> ), .B(n448), .C(\readoutR0<4> ), .D(n449), 
        .Y(n48) );
  NAND3X1 U89 ( .A(n393), .B(n425), .C(n55), .Y(n480) );
  AOI22X1 U90 ( .A(\readoutR7<3> ), .B(n9), .C(\readoutR6<3> ), .D(n8), .Y(n57) );
  AOI22X1 U91 ( .A(\readoutR5<3> ), .B(n11), .C(\readoutR4<3> ), .D(n10), .Y(
        n56) );
  AOI22X1 U92 ( .A(\readoutR3<3> ), .B(n450), .C(\readoutR2<3> ), .D(n451), 
        .Y(n54) );
  AOI22X1 U93 ( .A(\readoutR1<3> ), .B(n448), .C(\readoutR0<3> ), .D(n449), 
        .Y(n53) );
  NAND3X1 U94 ( .A(n392), .B(n424), .C(n60), .Y(n481) );
  AOI22X1 U95 ( .A(\readoutR7<2> ), .B(n9), .C(\readoutR6<2> ), .D(n8), .Y(n62) );
  AOI22X1 U96 ( .A(\readoutR5<2> ), .B(n11), .C(\readoutR4<2> ), .D(n10), .Y(
        n61) );
  AOI22X1 U97 ( .A(\readoutR3<2> ), .B(n450), .C(\readoutR2<2> ), .D(n451), 
        .Y(n59) );
  AOI22X1 U98 ( .A(\readoutR1<2> ), .B(n448), .C(\readoutR0<2> ), .D(n449), 
        .Y(n58) );
  NAND3X1 U99 ( .A(n391), .B(n423), .C(n65), .Y(n482) );
  AOI22X1 U100 ( .A(\readoutR7<1> ), .B(n9), .C(\readoutR6<1> ), .D(n8), .Y(
        n67) );
  AOI22X1 U101 ( .A(\readoutR5<1> ), .B(n11), .C(\readoutR4<1> ), .D(n10), .Y(
        n66) );
  AOI22X1 U102 ( .A(\readoutR3<1> ), .B(n450), .C(\readoutR2<1> ), .D(n451), 
        .Y(n64) );
  AOI22X1 U103 ( .A(\readoutR1<1> ), .B(n448), .C(\readoutR0<1> ), .D(n449), 
        .Y(n63) );
  NAND3X1 U104 ( .A(n390), .B(n422), .C(n70), .Y(n468) );
  AOI22X1 U105 ( .A(\readoutR7<15> ), .B(n9), .C(\readoutR6<15> ), .D(n8), .Y(
        n72) );
  AOI22X1 U106 ( .A(\readoutR5<15> ), .B(n11), .C(\readoutR4<15> ), .D(n10), 
        .Y(n71) );
  AOI22X1 U107 ( .A(\readoutR3<15> ), .B(n450), .C(\readoutR2<15> ), .D(n451), 
        .Y(n69) );
  AOI22X1 U108 ( .A(\readoutR1<15> ), .B(n448), .C(\readoutR0<15> ), .D(n449), 
        .Y(n68) );
  NAND3X1 U109 ( .A(n389), .B(n421), .C(n75), .Y(n469) );
  AOI22X1 U110 ( .A(\readoutR7<14> ), .B(n9), .C(\readoutR6<14> ), .D(n8), .Y(
        n77) );
  AOI22X1 U111 ( .A(\readoutR5<14> ), .B(n11), .C(\readoutR4<14> ), .D(n10), 
        .Y(n76) );
  AOI22X1 U112 ( .A(\readoutR3<14> ), .B(n450), .C(\readoutR2<14> ), .D(n451), 
        .Y(n74) );
  AOI22X1 U113 ( .A(\readoutR1<14> ), .B(n448), .C(\readoutR0<14> ), .D(n449), 
        .Y(n73) );
  NAND3X1 U114 ( .A(n388), .B(n420), .C(n80), .Y(n470) );
  AOI22X1 U115 ( .A(\readoutR7<13> ), .B(n9), .C(\readoutR6<13> ), .D(n8), .Y(
        n82) );
  AOI22X1 U116 ( .A(\readoutR5<13> ), .B(n11), .C(\readoutR4<13> ), .D(n10), 
        .Y(n81) );
  AOI22X1 U117 ( .A(\readoutR3<13> ), .B(n450), .C(\readoutR2<13> ), .D(n451), 
        .Y(n79) );
  AOI22X1 U118 ( .A(\readoutR1<13> ), .B(n448), .C(\readoutR0<13> ), .D(n449), 
        .Y(n78) );
  NAND3X1 U119 ( .A(n387), .B(n419), .C(n85), .Y(n471) );
  AOI22X1 U120 ( .A(\readoutR7<12> ), .B(n9), .C(\readoutR6<12> ), .D(n8), .Y(
        n87) );
  AOI22X1 U121 ( .A(\readoutR5<12> ), .B(n11), .C(\readoutR4<12> ), .D(n10), 
        .Y(n86) );
  AOI22X1 U122 ( .A(\readoutR3<12> ), .B(n450), .C(\readoutR2<12> ), .D(n451), 
        .Y(n84) );
  AOI22X1 U123 ( .A(\readoutR1<12> ), .B(n448), .C(\readoutR0<12> ), .D(n449), 
        .Y(n83) );
  NAND3X1 U124 ( .A(n386), .B(n418), .C(n90), .Y(n472) );
  AOI22X1 U125 ( .A(\readoutR7<11> ), .B(n9), .C(\readoutR6<11> ), .D(n8), .Y(
        n92) );
  AOI22X1 U126 ( .A(\readoutR5<11> ), .B(n11), .C(\readoutR4<11> ), .D(n10), 
        .Y(n91) );
  AOI22X1 U127 ( .A(\readoutR3<11> ), .B(n450), .C(\readoutR2<11> ), .D(n451), 
        .Y(n89) );
  AOI22X1 U128 ( .A(\readoutR1<11> ), .B(n448), .C(\readoutR0<11> ), .D(n449), 
        .Y(n88) );
  NAND3X1 U129 ( .A(n385), .B(n417), .C(n95), .Y(n473) );
  AOI22X1 U130 ( .A(\readoutR7<10> ), .B(n9), .C(\readoutR6<10> ), .D(n8), .Y(
        n97) );
  AOI22X1 U131 ( .A(\readoutR5<10> ), .B(n11), .C(\readoutR4<10> ), .D(n10), 
        .Y(n96) );
  AOI22X1 U132 ( .A(\readoutR3<10> ), .B(n450), .C(\readoutR2<10> ), .D(n451), 
        .Y(n94) );
  AOI22X1 U133 ( .A(\readoutR1<10> ), .B(n448), .C(\readoutR0<10> ), .D(n449), 
        .Y(n93) );
  NAND3X1 U134 ( .A(n384), .B(n416), .C(n100), .Y(n483) );
  AOI22X1 U135 ( .A(\readoutR7<0> ), .B(n9), .C(\readoutR6<0> ), .D(n8), .Y(
        n102) );
  NAND3X1 U136 ( .A(\read2regsel<1> ), .B(n13), .C(\read2regsel<2> ), .Y(n103)
         );
  NAND3X1 U137 ( .A(\read2regsel<1> ), .B(\read2regsel<0> ), .C(
        \read2regsel<2> ), .Y(n104) );
  AOI22X1 U138 ( .A(\readoutR5<0> ), .B(n11), .C(\readoutR4<0> ), .D(n10), .Y(
        n101) );
  NAND3X1 U139 ( .A(n13), .B(n12), .C(\read2regsel<2> ), .Y(n105) );
  NAND3X1 U140 ( .A(\read2regsel<0> ), .B(n12), .C(\read2regsel<2> ), .Y(n106)
         );
  AOI22X1 U141 ( .A(\readoutR3<0> ), .B(n450), .C(\readoutR2<0> ), .D(n451), 
        .Y(n99) );
  NOR3X1 U142 ( .A(\read2regsel<0> ), .B(\read2regsel<2> ), .C(n12), .Y(n25)
         );
  NOR3X1 U143 ( .A(n13), .B(\read2regsel<2> ), .C(n12), .Y(n24) );
  AOI22X1 U144 ( .A(\readoutR1<0> ), .B(n448), .C(\readoutR0<0> ), .D(n449), 
        .Y(n98) );
  NOR3X1 U145 ( .A(\read2regsel<1> ), .B(\read2regsel<2> ), .C(
        \read2regsel<0> ), .Y(n27) );
  NOR3X1 U146 ( .A(\read2regsel<1> ), .B(\read2regsel<2> ), .C(n13), .Y(n26)
         );
  NAND3X1 U147 ( .A(n383), .B(n415), .C(n109), .Y(n458) );
  AOI22X1 U148 ( .A(n3), .B(\readoutR7<9> ), .C(n2), .D(\readoutR6<9> ), .Y(
        n111) );
  AOI22X1 U149 ( .A(n5), .B(\readoutR5<9> ), .C(n4), .D(\readoutR4<9> ), .Y(
        n110) );
  AOI22X1 U150 ( .A(n446), .B(\readoutR3<9> ), .C(n447), .D(\readoutR2<9> ), 
        .Y(n108) );
  AOI22X1 U151 ( .A(n444), .B(\readoutR1<9> ), .C(n445), .D(\readoutR0<9> ), 
        .Y(n107) );
  NAND3X1 U152 ( .A(n382), .B(n414), .C(n118), .Y(n459) );
  AOI22X1 U153 ( .A(n3), .B(\readoutR7<8> ), .C(n2), .D(\readoutR6<8> ), .Y(
        n120) );
  AOI22X1 U154 ( .A(n5), .B(\readoutR5<8> ), .C(n4), .D(\readoutR4<8> ), .Y(
        n119) );
  AOI22X1 U155 ( .A(n446), .B(\readoutR3<8> ), .C(n447), .D(\readoutR2<8> ), 
        .Y(n117) );
  AOI22X1 U156 ( .A(n444), .B(\readoutR1<8> ), .C(n445), .D(\readoutR0<8> ), 
        .Y(n116) );
  NAND3X1 U157 ( .A(n381), .B(n413), .C(n123), .Y(n460) );
  AOI22X1 U158 ( .A(n3), .B(\readoutR7<7> ), .C(n2), .D(\readoutR6<7> ), .Y(
        n125) );
  AOI22X1 U159 ( .A(n5), .B(\readoutR5<7> ), .C(n4), .D(\readoutR4<7> ), .Y(
        n124) );
  AOI22X1 U160 ( .A(n446), .B(\readoutR3<7> ), .C(n447), .D(\readoutR2<7> ), 
        .Y(n122) );
  AOI22X1 U161 ( .A(n444), .B(\readoutR1<7> ), .C(n445), .D(\readoutR0<7> ), 
        .Y(n121) );
  NAND3X1 U162 ( .A(n380), .B(n412), .C(n128), .Y(n461) );
  AOI22X1 U163 ( .A(n3), .B(\readoutR7<6> ), .C(n2), .D(\readoutR6<6> ), .Y(
        n130) );
  AOI22X1 U164 ( .A(n5), .B(\readoutR5<6> ), .C(n4), .D(\readoutR4<6> ), .Y(
        n129) );
  AOI22X1 U165 ( .A(n446), .B(\readoutR3<6> ), .C(n447), .D(\readoutR2<6> ), 
        .Y(n127) );
  AOI22X1 U166 ( .A(n444), .B(\readoutR1<6> ), .C(n445), .D(\readoutR0<6> ), 
        .Y(n126) );
  NAND3X1 U167 ( .A(n379), .B(n411), .C(n133), .Y(n462) );
  AOI22X1 U168 ( .A(n3), .B(\readoutR7<5> ), .C(n2), .D(\readoutR6<5> ), .Y(
        n135) );
  AOI22X1 U169 ( .A(n5), .B(\readoutR5<5> ), .C(n4), .D(\readoutR4<5> ), .Y(
        n134) );
  AOI22X1 U170 ( .A(n446), .B(\readoutR3<5> ), .C(n447), .D(\readoutR2<5> ), 
        .Y(n132) );
  AOI22X1 U171 ( .A(n444), .B(\readoutR1<5> ), .C(n445), .D(\readoutR0<5> ), 
        .Y(n131) );
  NAND3X1 U172 ( .A(n378), .B(n410), .C(n138), .Y(n463) );
  AOI22X1 U173 ( .A(n3), .B(\readoutR7<4> ), .C(n2), .D(\readoutR6<4> ), .Y(
        n140) );
  AOI22X1 U174 ( .A(n5), .B(\readoutR5<4> ), .C(n4), .D(\readoutR4<4> ), .Y(
        n139) );
  AOI22X1 U175 ( .A(n446), .B(\readoutR3<4> ), .C(n447), .D(\readoutR2<4> ), 
        .Y(n137) );
  AOI22X1 U176 ( .A(n444), .B(\readoutR1<4> ), .C(n445), .D(\readoutR0<4> ), 
        .Y(n136) );
  NAND3X1 U177 ( .A(n377), .B(n409), .C(n143), .Y(n464) );
  AOI22X1 U178 ( .A(n3), .B(\readoutR7<3> ), .C(n2), .D(\readoutR6<3> ), .Y(
        n145) );
  AOI22X1 U179 ( .A(n5), .B(\readoutR5<3> ), .C(n4), .D(\readoutR4<3> ), .Y(
        n144) );
  AOI22X1 U180 ( .A(n446), .B(\readoutR3<3> ), .C(n447), .D(\readoutR2<3> ), 
        .Y(n142) );
  AOI22X1 U181 ( .A(n444), .B(\readoutR1<3> ), .C(n445), .D(\readoutR0<3> ), 
        .Y(n141) );
  NAND3X1 U182 ( .A(n376), .B(n408), .C(n148), .Y(n465) );
  AOI22X1 U183 ( .A(n3), .B(\readoutR7<2> ), .C(n2), .D(\readoutR6<2> ), .Y(
        n150) );
  AOI22X1 U184 ( .A(n5), .B(\readoutR5<2> ), .C(n4), .D(\readoutR4<2> ), .Y(
        n149) );
  AOI22X1 U185 ( .A(n446), .B(\readoutR3<2> ), .C(n447), .D(\readoutR2<2> ), 
        .Y(n147) );
  AOI22X1 U186 ( .A(n444), .B(\readoutR1<2> ), .C(n445), .D(\readoutR0<2> ), 
        .Y(n146) );
  NAND3X1 U187 ( .A(n375), .B(n407), .C(n153), .Y(n466) );
  AOI22X1 U188 ( .A(n3), .B(\readoutR7<1> ), .C(n2), .D(\readoutR6<1> ), .Y(
        n155) );
  AOI22X1 U189 ( .A(n5), .B(\readoutR5<1> ), .C(n4), .D(\readoutR4<1> ), .Y(
        n154) );
  AOI22X1 U190 ( .A(n446), .B(\readoutR3<1> ), .C(n447), .D(\readoutR2<1> ), 
        .Y(n152) );
  AOI22X1 U191 ( .A(n444), .B(\readoutR1<1> ), .C(n445), .D(\readoutR0<1> ), 
        .Y(n151) );
  NAND3X1 U192 ( .A(n374), .B(n406), .C(n158), .Y(n452) );
  AOI22X1 U193 ( .A(n3), .B(\readoutR7<15> ), .C(n2), .D(\readoutR6<15> ), .Y(
        n160) );
  AOI22X1 U194 ( .A(n5), .B(\readoutR5<15> ), .C(n4), .D(\readoutR4<15> ), .Y(
        n159) );
  AOI22X1 U195 ( .A(n446), .B(\readoutR3<15> ), .C(n447), .D(\readoutR2<15> ), 
        .Y(n157) );
  AOI22X1 U196 ( .A(n444), .B(\readoutR1<15> ), .C(n445), .D(\readoutR0<15> ), 
        .Y(n156) );
  NAND3X1 U197 ( .A(n373), .B(n405), .C(n163), .Y(n453) );
  AOI22X1 U198 ( .A(n3), .B(\readoutR7<14> ), .C(n2), .D(\readoutR6<14> ), .Y(
        n165) );
  AOI22X1 U199 ( .A(n5), .B(\readoutR5<14> ), .C(n4), .D(\readoutR4<14> ), .Y(
        n164) );
  AOI22X1 U200 ( .A(n446), .B(\readoutR3<14> ), .C(n447), .D(\readoutR2<14> ), 
        .Y(n162) );
  AOI22X1 U201 ( .A(n444), .B(\readoutR1<14> ), .C(n445), .D(\readoutR0<14> ), 
        .Y(n161) );
  NAND3X1 U202 ( .A(n372), .B(n404), .C(n168), .Y(n454) );
  AOI22X1 U203 ( .A(n3), .B(\readoutR7<13> ), .C(n2), .D(\readoutR6<13> ), .Y(
        n170) );
  AOI22X1 U204 ( .A(n5), .B(\readoutR5<13> ), .C(n4), .D(\readoutR4<13> ), .Y(
        n169) );
  AOI22X1 U205 ( .A(n446), .B(\readoutR3<13> ), .C(n447), .D(\readoutR2<13> ), 
        .Y(n167) );
  AOI22X1 U206 ( .A(n444), .B(\readoutR1<13> ), .C(n445), .D(\readoutR0<13> ), 
        .Y(n166) );
  NAND3X1 U207 ( .A(n371), .B(n403), .C(n173), .Y(n455) );
  AOI22X1 U208 ( .A(n3), .B(\readoutR7<12> ), .C(n2), .D(\readoutR6<12> ), .Y(
        n175) );
  AOI22X1 U209 ( .A(n5), .B(\readoutR5<12> ), .C(n4), .D(\readoutR4<12> ), .Y(
        n174) );
  AOI22X1 U210 ( .A(n446), .B(\readoutR3<12> ), .C(n447), .D(\readoutR2<12> ), 
        .Y(n172) );
  AOI22X1 U211 ( .A(n444), .B(\readoutR1<12> ), .C(n445), .D(\readoutR0<12> ), 
        .Y(n171) );
  NAND3X1 U212 ( .A(n370), .B(n402), .C(n178), .Y(n456) );
  AOI22X1 U213 ( .A(n3), .B(\readoutR7<11> ), .C(n2), .D(\readoutR6<11> ), .Y(
        n180) );
  AOI22X1 U214 ( .A(n5), .B(\readoutR5<11> ), .C(n4), .D(\readoutR4<11> ), .Y(
        n179) );
  AOI22X1 U215 ( .A(n446), .B(\readoutR3<11> ), .C(n447), .D(\readoutR2<11> ), 
        .Y(n177) );
  AOI22X1 U216 ( .A(n444), .B(\readoutR1<11> ), .C(n445), .D(\readoutR0<11> ), 
        .Y(n176) );
  NAND3X1 U217 ( .A(n369), .B(n401), .C(n183), .Y(n457) );
  AOI22X1 U218 ( .A(n3), .B(\readoutR7<10> ), .C(n2), .D(\readoutR6<10> ), .Y(
        n185) );
  AOI22X1 U219 ( .A(n5), .B(\readoutR5<10> ), .C(n4), .D(\readoutR4<10> ), .Y(
        n184) );
  AOI22X1 U220 ( .A(n446), .B(\readoutR3<10> ), .C(n447), .D(\readoutR2<10> ), 
        .Y(n182) );
  AOI22X1 U221 ( .A(n444), .B(\readoutR1<10> ), .C(n445), .D(\readoutR0<10> ), 
        .Y(n181) );
  NAND3X1 U222 ( .A(n368), .B(n400), .C(n188), .Y(n467) );
  AOI22X1 U223 ( .A(n3), .B(\readoutR7<0> ), .C(n2), .D(\readoutR6<0> ), .Y(
        n190) );
  NAND3X1 U224 ( .A(\read1regsel<1> ), .B(n7), .C(\read1regsel<2> ), .Y(n191)
         );
  NAND3X1 U225 ( .A(\read1regsel<1> ), .B(\read1regsel<0> ), .C(
        \read1regsel<2> ), .Y(n192) );
  AOI22X1 U226 ( .A(n5), .B(\readoutR5<0> ), .C(n4), .D(\readoutR4<0> ), .Y(
        n189) );
  NAND3X1 U227 ( .A(n7), .B(n6), .C(\read1regsel<2> ), .Y(n193) );
  NAND3X1 U228 ( .A(\read1regsel<0> ), .B(n6), .C(\read1regsel<2> ), .Y(n194)
         );
  AOI22X1 U229 ( .A(n446), .B(\readoutR3<0> ), .C(n447), .D(\readoutR2<0> ), 
        .Y(n187) );
  NOR3X1 U230 ( .A(\read1regsel<0> ), .B(\read1regsel<2> ), .C(n6), .Y(n113)
         );
  NOR3X1 U231 ( .A(n7), .B(\read1regsel<2> ), .C(n6), .Y(n112) );
  AOI22X1 U232 ( .A(n444), .B(\readoutR1<0> ), .C(n445), .D(\readoutR0<0> ), 
        .Y(n186) );
  NOR3X1 U233 ( .A(\read1regsel<1> ), .B(\read1regsel<2> ), .C(
        \read1regsel<0> ), .Y(n115) );
  NOR3X1 U234 ( .A(\read1regsel<1> ), .B(\read1regsel<2> ), .C(n7), .Y(n114)
         );
  BUFX2 U18 ( .A(n115), .Y(n445) );
  BUFX2 U19 ( .A(n113), .Y(n447) );
  BUFX2 U20 ( .A(n27), .Y(n449) );
  BUFX2 U21 ( .A(n25), .Y(n451) );
  AND2X1 U22 ( .A(write), .B(n16), .Y(n440) );
  INVX1 U23 ( .A(\writeregsel<0> ), .Y(n16) );
  AND2X1 U24 ( .A(\writeregsel<0> ), .B(write), .Y(n442) );
  INVX1 U25 ( .A(\writeregsel<2> ), .Y(n14) );
  INVX1 U26 ( .A(\writeregsel<1> ), .Y(n15) );
  INVX1 U27 ( .A(\read2regsel<1> ), .Y(n12) );
  AND2X1 U28 ( .A(n17), .B(n273), .Y(n188) );
  AND2X1 U29 ( .A(n195), .B(n275), .Y(n183) );
  AND2X1 U30 ( .A(n197), .B(n277), .Y(n178) );
  AND2X1 U31 ( .A(n199), .B(n279), .Y(n173) );
  AND2X1 U32 ( .A(n201), .B(n281), .Y(n168) );
  AND2X1 U33 ( .A(n203), .B(n283), .Y(n163) );
  AND2X1 U34 ( .A(n205), .B(n285), .Y(n158) );
  AND2X1 U35 ( .A(n207), .B(n287), .Y(n153) );
  AND2X1 U36 ( .A(n209), .B(n289), .Y(n148) );
  AND2X1 U37 ( .A(n211), .B(n291), .Y(n143) );
  AND2X1 U40 ( .A(n213), .B(n293), .Y(n138) );
  AND2X1 U41 ( .A(n215), .B(n295), .Y(n133) );
  AND2X1 U42 ( .A(n217), .B(n297), .Y(n128) );
  AND2X1 U43 ( .A(n219), .B(n299), .Y(n123) );
  AND2X1 U44 ( .A(n221), .B(n301), .Y(n118) );
  AND2X1 U46 ( .A(n223), .B(n303), .Y(n109) );
  INVX1 U47 ( .A(n189), .Y(n1) );
  INVX1 U48 ( .A(n1), .Y(n17) );
  INVX1 U56 ( .A(n184), .Y(n18) );
  INVX1 U58 ( .A(n18), .Y(n195) );
  INVX1 U235 ( .A(n179), .Y(n196) );
  INVX1 U236 ( .A(n196), .Y(n197) );
  INVX1 U237 ( .A(n174), .Y(n198) );
  INVX1 U238 ( .A(n198), .Y(n199) );
  INVX1 U239 ( .A(n169), .Y(n200) );
  INVX1 U240 ( .A(n200), .Y(n201) );
  INVX1 U241 ( .A(n164), .Y(n202) );
  INVX1 U242 ( .A(n202), .Y(n203) );
  INVX1 U243 ( .A(n159), .Y(n204) );
  INVX1 U244 ( .A(n204), .Y(n205) );
  INVX1 U245 ( .A(n154), .Y(n206) );
  INVX1 U246 ( .A(n206), .Y(n207) );
  INVX1 U247 ( .A(n149), .Y(n208) );
  INVX1 U248 ( .A(n208), .Y(n209) );
  INVX1 U249 ( .A(n144), .Y(n210) );
  INVX1 U250 ( .A(n210), .Y(n211) );
  INVX1 U251 ( .A(n139), .Y(n212) );
  INVX1 U252 ( .A(n212), .Y(n213) );
  INVX1 U253 ( .A(n134), .Y(n214) );
  INVX1 U254 ( .A(n214), .Y(n215) );
  INVX1 U255 ( .A(n129), .Y(n216) );
  INVX1 U256 ( .A(n216), .Y(n217) );
  INVX1 U257 ( .A(n124), .Y(n218) );
  INVX1 U258 ( .A(n218), .Y(n219) );
  INVX1 U259 ( .A(n119), .Y(n220) );
  INVX1 U260 ( .A(n220), .Y(n221) );
  INVX1 U261 ( .A(n110), .Y(n222) );
  INVX1 U262 ( .A(n222), .Y(n223) );
  INVX1 U263 ( .A(n101), .Y(n224) );
  INVX1 U264 ( .A(n224), .Y(n225) );
  INVX1 U265 ( .A(n96), .Y(n226) );
  INVX1 U266 ( .A(n226), .Y(n227) );
  INVX1 U267 ( .A(n91), .Y(n228) );
  INVX1 U268 ( .A(n228), .Y(n229) );
  INVX1 U269 ( .A(n86), .Y(n230) );
  INVX1 U270 ( .A(n230), .Y(n231) );
  INVX1 U271 ( .A(n81), .Y(n232) );
  INVX1 U272 ( .A(n232), .Y(n233) );
  INVX1 U273 ( .A(n76), .Y(n234) );
  INVX1 U274 ( .A(n234), .Y(n235) );
  INVX1 U275 ( .A(n71), .Y(n236) );
  INVX1 U276 ( .A(n236), .Y(n237) );
  INVX1 U277 ( .A(n66), .Y(n238) );
  INVX1 U278 ( .A(n238), .Y(n239) );
  INVX1 U279 ( .A(n61), .Y(n240) );
  INVX1 U280 ( .A(n240), .Y(n241) );
  INVX1 U281 ( .A(n56), .Y(n242) );
  INVX1 U282 ( .A(n242), .Y(n243) );
  INVX1 U283 ( .A(n51), .Y(n244) );
  INVX1 U284 ( .A(n244), .Y(n245) );
  INVX1 U285 ( .A(n46), .Y(n246) );
  INVX1 U286 ( .A(n246), .Y(n247) );
  INVX1 U287 ( .A(n41), .Y(n248) );
  INVX1 U288 ( .A(n248), .Y(n249) );
  INVX1 U289 ( .A(n36), .Y(n250) );
  INVX1 U290 ( .A(n250), .Y(n251) );
  INVX1 U291 ( .A(n31), .Y(n252) );
  INVX1 U292 ( .A(n252), .Y(n253) );
  INVX1 U293 ( .A(n22), .Y(n254) );
  INVX1 U294 ( .A(n254), .Y(n255) );
  BUFX2 U295 ( .A(n102), .Y(n256) );
  BUFX2 U296 ( .A(n97), .Y(n257) );
  BUFX2 U297 ( .A(n92), .Y(n258) );
  BUFX2 U298 ( .A(n87), .Y(n259) );
  BUFX2 U299 ( .A(n82), .Y(n260) );
  BUFX2 U300 ( .A(n77), .Y(n261) );
  BUFX2 U301 ( .A(n72), .Y(n262) );
  BUFX2 U302 ( .A(n67), .Y(n263) );
  BUFX2 U303 ( .A(n62), .Y(n264) );
  BUFX2 U304 ( .A(n57), .Y(n265) );
  BUFX2 U305 ( .A(n52), .Y(n266) );
  BUFX2 U306 ( .A(n47), .Y(n267) );
  BUFX2 U307 ( .A(n42), .Y(n268) );
  BUFX2 U308 ( .A(n37), .Y(n269) );
  BUFX2 U309 ( .A(n32), .Y(n270) );
  BUFX2 U310 ( .A(n23), .Y(n271) );
  BUFX2 U311 ( .A(n114), .Y(n444) );
  BUFX2 U312 ( .A(n112), .Y(n446) );
  BUFX2 U313 ( .A(n26), .Y(n448) );
  BUFX2 U314 ( .A(n24), .Y(n450) );
  INVX1 U315 ( .A(n190), .Y(n272) );
  INVX1 U316 ( .A(n272), .Y(n273) );
  INVX1 U317 ( .A(n185), .Y(n274) );
  INVX1 U318 ( .A(n274), .Y(n275) );
  INVX1 U319 ( .A(n180), .Y(n276) );
  INVX1 U320 ( .A(n276), .Y(n277) );
  INVX1 U321 ( .A(n175), .Y(n278) );
  INVX1 U322 ( .A(n278), .Y(n279) );
  INVX1 U323 ( .A(n170), .Y(n280) );
  INVX1 U324 ( .A(n280), .Y(n281) );
  INVX1 U325 ( .A(n165), .Y(n282) );
  INVX1 U326 ( .A(n282), .Y(n283) );
  INVX1 U327 ( .A(n160), .Y(n284) );
  INVX1 U328 ( .A(n284), .Y(n285) );
  INVX1 U329 ( .A(n155), .Y(n286) );
  INVX1 U330 ( .A(n286), .Y(n287) );
  INVX1 U331 ( .A(n150), .Y(n288) );
  INVX1 U332 ( .A(n288), .Y(n289) );
  INVX1 U333 ( .A(n145), .Y(n290) );
  INVX1 U334 ( .A(n290), .Y(n291) );
  INVX1 U335 ( .A(n140), .Y(n292) );
  INVX1 U336 ( .A(n292), .Y(n293) );
  INVX1 U337 ( .A(n135), .Y(n294) );
  INVX1 U338 ( .A(n294), .Y(n295) );
  INVX1 U339 ( .A(n130), .Y(n296) );
  INVX1 U340 ( .A(n296), .Y(n297) );
  INVX1 U341 ( .A(n125), .Y(n298) );
  INVX1 U342 ( .A(n298), .Y(n299) );
  INVX1 U343 ( .A(n120), .Y(n300) );
  INVX1 U344 ( .A(n300), .Y(n301) );
  INVX1 U345 ( .A(n111), .Y(n302) );
  INVX1 U346 ( .A(n302), .Y(n303) );
  INVX1 U347 ( .A(n467), .Y(n304) );
  INVX1 U348 ( .A(n304), .Y(\read1data<0> ) );
  INVX1 U349 ( .A(n457), .Y(n306) );
  INVX1 U350 ( .A(n306), .Y(\read1data<10> ) );
  INVX1 U351 ( .A(n456), .Y(n308) );
  INVX1 U352 ( .A(n308), .Y(\read1data<11> ) );
  INVX1 U353 ( .A(n455), .Y(n310) );
  INVX1 U354 ( .A(n310), .Y(\read1data<12> ) );
  INVX1 U355 ( .A(n454), .Y(n312) );
  INVX1 U356 ( .A(n312), .Y(\read1data<13> ) );
  INVX1 U357 ( .A(n453), .Y(n314) );
  INVX1 U358 ( .A(n314), .Y(\read1data<14> ) );
  INVX1 U359 ( .A(n452), .Y(n316) );
  INVX1 U360 ( .A(n316), .Y(\read1data<15> ) );
  INVX1 U361 ( .A(n466), .Y(n318) );
  INVX1 U362 ( .A(n318), .Y(\read1data<1> ) );
  INVX1 U363 ( .A(n465), .Y(n320) );
  INVX1 U364 ( .A(n320), .Y(\read1data<2> ) );
  INVX1 U365 ( .A(n464), .Y(n322) );
  INVX1 U366 ( .A(n322), .Y(\read1data<3> ) );
  INVX1 U367 ( .A(n463), .Y(n324) );
  INVX1 U368 ( .A(n324), .Y(\read1data<4> ) );
  INVX1 U369 ( .A(n462), .Y(n326) );
  INVX1 U370 ( .A(n326), .Y(\read1data<5> ) );
  INVX1 U371 ( .A(n461), .Y(n328) );
  INVX1 U372 ( .A(n328), .Y(\read1data<6> ) );
  INVX1 U373 ( .A(n460), .Y(n330) );
  INVX1 U374 ( .A(n330), .Y(\read1data<7> ) );
  INVX1 U375 ( .A(n459), .Y(n332) );
  INVX1 U376 ( .A(n332), .Y(\read1data<8> ) );
  INVX1 U377 ( .A(n458), .Y(n334) );
  INVX1 U378 ( .A(n334), .Y(\read1data<9> ) );
  INVX1 U379 ( .A(n483), .Y(n336) );
  INVX1 U380 ( .A(n336), .Y(\read2data<0> ) );
  INVX1 U381 ( .A(n473), .Y(n338) );
  INVX1 U382 ( .A(n338), .Y(\read2data<10> ) );
  INVX1 U383 ( .A(n472), .Y(n340) );
  INVX1 U384 ( .A(n340), .Y(\read2data<11> ) );
  INVX1 U385 ( .A(n471), .Y(n342) );
  INVX1 U386 ( .A(n342), .Y(\read2data<12> ) );
  INVX1 U387 ( .A(n470), .Y(n344) );
  INVX1 U388 ( .A(n344), .Y(\read2data<13> ) );
  INVX1 U389 ( .A(n469), .Y(n346) );
  INVX1 U390 ( .A(n346), .Y(\read2data<14> ) );
  INVX1 U391 ( .A(n468), .Y(n348) );
  INVX1 U392 ( .A(n348), .Y(\read2data<15> ) );
  INVX1 U393 ( .A(n482), .Y(n350) );
  INVX1 U394 ( .A(n350), .Y(\read2data<1> ) );
  INVX1 U395 ( .A(n481), .Y(n352) );
  INVX1 U396 ( .A(n352), .Y(\read2data<2> ) );
  INVX1 U397 ( .A(n480), .Y(n354) );
  INVX1 U398 ( .A(n354), .Y(\read2data<3> ) );
  INVX1 U399 ( .A(n479), .Y(n356) );
  INVX1 U400 ( .A(n356), .Y(\read2data<4> ) );
  INVX1 U401 ( .A(n478), .Y(n358) );
  INVX1 U402 ( .A(n358), .Y(\read2data<5> ) );
  INVX1 U403 ( .A(n477), .Y(n360) );
  INVX1 U404 ( .A(n360), .Y(\read2data<6> ) );
  INVX1 U405 ( .A(n476), .Y(n362) );
  INVX1 U406 ( .A(n362), .Y(\read2data<7> ) );
  INVX1 U407 ( .A(n475), .Y(n364) );
  INVX1 U408 ( .A(n364), .Y(\read2data<8> ) );
  INVX1 U409 ( .A(n474), .Y(n366) );
  INVX1 U410 ( .A(n366), .Y(\read2data<9> ) );
  BUFX2 U411 ( .A(n186), .Y(n368) );
  BUFX2 U412 ( .A(n181), .Y(n369) );
  BUFX2 U413 ( .A(n176), .Y(n370) );
  BUFX2 U414 ( .A(n171), .Y(n371) );
  BUFX2 U415 ( .A(n166), .Y(n372) );
  BUFX2 U416 ( .A(n161), .Y(n373) );
  BUFX2 U417 ( .A(n156), .Y(n374) );
  BUFX2 U418 ( .A(n151), .Y(n375) );
  BUFX2 U419 ( .A(n146), .Y(n376) );
  BUFX2 U420 ( .A(n141), .Y(n377) );
  BUFX2 U421 ( .A(n136), .Y(n378) );
  BUFX2 U422 ( .A(n131), .Y(n379) );
  BUFX2 U423 ( .A(n126), .Y(n380) );
  BUFX2 U424 ( .A(n121), .Y(n381) );
  BUFX2 U425 ( .A(n116), .Y(n382) );
  BUFX2 U426 ( .A(n107), .Y(n383) );
  BUFX2 U427 ( .A(n98), .Y(n384) );
  BUFX2 U428 ( .A(n93), .Y(n385) );
  BUFX2 U429 ( .A(n88), .Y(n386) );
  BUFX2 U430 ( .A(n83), .Y(n387) );
  BUFX2 U431 ( .A(n78), .Y(n388) );
  BUFX2 U432 ( .A(n73), .Y(n389) );
  BUFX2 U433 ( .A(n68), .Y(n390) );
  BUFX2 U434 ( .A(n63), .Y(n391) );
  BUFX2 U435 ( .A(n58), .Y(n392) );
  BUFX2 U436 ( .A(n53), .Y(n393) );
  BUFX2 U437 ( .A(n48), .Y(n394) );
  BUFX2 U438 ( .A(n43), .Y(n395) );
  BUFX2 U439 ( .A(n38), .Y(n396) );
  BUFX2 U440 ( .A(n33), .Y(n397) );
  BUFX2 U441 ( .A(n28), .Y(n398) );
  BUFX2 U442 ( .A(n19), .Y(n399) );
  BUFX2 U443 ( .A(n187), .Y(n400) );
  BUFX2 U444 ( .A(n182), .Y(n401) );
  BUFX2 U445 ( .A(n177), .Y(n402) );
  BUFX2 U446 ( .A(n172), .Y(n403) );
  BUFX2 U447 ( .A(n167), .Y(n404) );
  BUFX2 U448 ( .A(n162), .Y(n405) );
  BUFX2 U449 ( .A(n157), .Y(n406) );
  BUFX2 U450 ( .A(n152), .Y(n407) );
  BUFX2 U451 ( .A(n147), .Y(n408) );
  BUFX2 U452 ( .A(n142), .Y(n409) );
  BUFX2 U453 ( .A(n137), .Y(n410) );
  BUFX2 U454 ( .A(n132), .Y(n411) );
  BUFX2 U455 ( .A(n127), .Y(n412) );
  BUFX2 U456 ( .A(n122), .Y(n413) );
  BUFX2 U457 ( .A(n117), .Y(n414) );
  BUFX2 U458 ( .A(n108), .Y(n415) );
  BUFX2 U459 ( .A(n99), .Y(n416) );
  BUFX2 U460 ( .A(n94), .Y(n417) );
  BUFX2 U461 ( .A(n89), .Y(n418) );
  BUFX2 U462 ( .A(n84), .Y(n419) );
  BUFX2 U463 ( .A(n79), .Y(n420) );
  BUFX2 U464 ( .A(n74), .Y(n421) );
  BUFX2 U465 ( .A(n69), .Y(n422) );
  BUFX2 U466 ( .A(n64), .Y(n423) );
  BUFX2 U467 ( .A(n59), .Y(n424) );
  BUFX2 U468 ( .A(n54), .Y(n425) );
  BUFX2 U469 ( .A(n49), .Y(n426) );
  BUFX2 U470 ( .A(n44), .Y(n427) );
  BUFX2 U471 ( .A(n39), .Y(n428) );
  BUFX2 U472 ( .A(n34), .Y(n429) );
  BUFX2 U473 ( .A(n29), .Y(n430) );
  BUFX2 U474 ( .A(n20), .Y(n431) );
  BUFX2 U475 ( .A(n194), .Y(n432) );
  INVX1 U476 ( .A(n432), .Y(n5) );
  BUFX2 U477 ( .A(n193), .Y(n433) );
  INVX1 U478 ( .A(n433), .Y(n4) );
  BUFX2 U479 ( .A(n192), .Y(n434) );
  INVX1 U480 ( .A(n434), .Y(n3) );
  BUFX2 U481 ( .A(n191), .Y(n435) );
  INVX1 U482 ( .A(n435), .Y(n2) );
  BUFX2 U483 ( .A(n106), .Y(n436) );
  INVX1 U484 ( .A(n436), .Y(n11) );
  BUFX2 U485 ( .A(n105), .Y(n437) );
  INVX1 U486 ( .A(n437), .Y(n10) );
  BUFX2 U487 ( .A(n104), .Y(n438) );
  INVX1 U488 ( .A(n438), .Y(n9) );
  BUFX2 U489 ( .A(n103), .Y(n439) );
  INVX1 U490 ( .A(n439), .Y(n8) );
  INVX1 U491 ( .A(n440), .Y(n441) );
  INVX1 U492 ( .A(n442), .Y(n443) );
endmodule


module dff_597 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_596 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_595 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_594 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_593 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_592 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_591 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_590 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_589 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_588 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_587 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_586 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_585 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_584 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_583 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_582 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_581 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_580 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_579 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_578 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_577 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_576 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_575 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_574 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_573 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_572 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_571 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_570 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_569 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_568 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_567 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_566 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_565 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_564 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_563 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_562 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_561 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_560 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_559 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_558 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_557 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_556 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_555 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_554 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_553 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_552 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_551 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_550 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_549 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_548 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_547 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_546 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_545 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_544 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_543 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_542 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_541 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_540 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_539 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_538 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_537 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_536 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_535 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_534 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_533 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_532 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_531 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_530 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_529 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_528 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_527 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_526 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_525 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_524 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_523 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_522 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_521 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_520 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_519 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_518 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_517 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_516 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_515 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_514 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_513 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_512 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_511 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_510 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_509 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_508 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_507 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_506 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_505 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_504 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_503 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_502 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_501 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_500 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_499 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_498 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_497 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_496 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_495 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_494 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_493 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_492 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_491 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_490 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_489 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_488 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_487 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_486 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_485 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_484 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_483 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_482 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_481 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_480 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_479 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_478 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_477 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_476 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_475 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_474 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_473 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_472 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_471 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_470 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_469 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_468 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_467 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_466 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_465 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_464 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_463 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_462 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_461 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_460 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_459 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_458 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_457 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_456 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_455 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_454 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_453 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_452 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module shifter ( .In({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), .Cnt({\Cnt<3> , \Cnt<2> , 
        \Cnt<1> , \Cnt<0> }), .Op({\Op<1> , \Op<0> }), .Out({\Out<15> , 
        \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> , \Out<9> , 
        \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , 
        \Out<1> , \Out<0> }) );
  input \In<15> , \In<14> , \In<13> , \In<12> , \In<11> , \In<10> , \In<9> ,
         \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , \In<3> , \In<2> ,
         \In<1> , \In<0> , \Cnt<3> , \Cnt<2> , \Cnt<1> , \Cnt<0> , \Op<1> ,
         \Op<0> ;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> ;
  wire   n772, n773, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n126, n128, n129, n130, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769;

  BUFX2 U2 ( .A(n186), .Y(n1) );
  INVX1 U3 ( .A(n92), .Y(n2) );
  INVX1 U4 ( .A(n2), .Y(n3) );
  INVX1 U5 ( .A(n538), .Y(n4) );
  INVX1 U6 ( .A(n130), .Y(n5) );
  INVX1 U7 ( .A(n170), .Y(n6) );
  INVX2 U8 ( .A(\Cnt<2> ), .Y(n66) );
  INVX1 U9 ( .A(n121), .Y(n584) );
  INVX1 U10 ( .A(n165), .Y(n7) );
  INVX1 U11 ( .A(n16), .Y(n8) );
  AND2X2 U12 ( .A(n293), .B(n447), .Y(n352) );
  INVX2 U13 ( .A(n138), .Y(n68) );
  AND2X2 U14 ( .A(\In<0> ), .B(n619), .Y(n9) );
  INVX1 U15 ( .A(n622), .Y(n26) );
  AND2X2 U16 ( .A(n214), .B(n205), .Y(n256) );
  INVX1 U17 ( .A(n682), .Y(n20) );
  INVX1 U18 ( .A(\In<1> ), .Y(n668) );
  AND2X1 U19 ( .A(n658), .B(n715), .Y(n175) );
  AND2X1 U20 ( .A(n193), .B(n561), .Y(n343) );
  INVX1 U21 ( .A(n83), .Y(n741) );
  INVX1 U22 ( .A(n556), .Y(n736) );
  OR2X1 U23 ( .A(n745), .B(n107), .Y(n57) );
  INVX4 U24 ( .A(n62), .Y(n763) );
  INVX1 U25 ( .A(n185), .Y(n10) );
  BUFX2 U26 ( .A(n68), .Y(n11) );
  INVX1 U27 ( .A(n576), .Y(n12) );
  INVX1 U28 ( .A(n100), .Y(n13) );
  INVX1 U29 ( .A(n152), .Y(n14) );
  INVX1 U30 ( .A(n372), .Y(n15) );
  OR2X1 U31 ( .A(n747), .B(n748), .Y(n372) );
  INVX1 U32 ( .A(n614), .Y(n16) );
  INVX1 U33 ( .A(n583), .Y(n17) );
  INVX1 U34 ( .A(n583), .Y(n582) );
  INVX1 U35 ( .A(n26), .Y(n18) );
  INVX1 U36 ( .A(n591), .Y(n19) );
  NOR3X1 U37 ( .A(n473), .B(n494), .C(n501), .Y(n21) );
  INVX1 U38 ( .A(n167), .Y(n22) );
  INVX1 U39 ( .A(n13), .Y(n23) );
  INVX1 U40 ( .A(n191), .Y(n24) );
  INVX1 U41 ( .A(n36), .Y(n25) );
  INVX1 U42 ( .A(n162), .Y(n27) );
  INVX1 U43 ( .A(n163), .Y(n28) );
  INVX1 U44 ( .A(n149), .Y(n29) );
  INVX1 U45 ( .A(n149), .Y(n585) );
  AND2X2 U46 ( .A(\In<1> ), .B(n619), .Y(n30) );
  INVX1 U47 ( .A(n105), .Y(n31) );
  AND2X2 U48 ( .A(n642), .B(n117), .Y(n32) );
  NOR2X1 U49 ( .A(n32), .B(n641), .Y(n643) );
  MUX2X1 U50 ( .B(n579), .A(n488), .S(n66), .Y(n735) );
  OR2X2 U51 ( .A(n212), .B(n34), .Y(n33) );
  INVX1 U52 ( .A(n33), .Y(n623) );
  INVX1 U53 ( .A(n673), .Y(n34) );
  AND2X1 U54 ( .A(n33), .B(n762), .Y(n334) );
  INVX1 U55 ( .A(n81), .Y(\Out<8> ) );
  BUFX2 U56 ( .A(n183), .Y(n35) );
  INVX1 U57 ( .A(n26), .Y(n36) );
  INVX1 U58 ( .A(n169), .Y(n37) );
  INVX1 U59 ( .A(n169), .Y(n38) );
  OR2X2 U60 ( .A(n116), .B(n160), .Y(n39) );
  INVX1 U61 ( .A(n113), .Y(n651) );
  AND2X2 U62 ( .A(n59), .B(n581), .Y(n40) );
  INVX1 U63 ( .A(n40), .Y(n46) );
  INVX1 U64 ( .A(n104), .Y(n41) );
  INVX1 U65 ( .A(n41), .Y(n42) );
  AND2X1 U66 ( .A(n463), .B(n64), .Y(n63) );
  INVX1 U67 ( .A(n756), .Y(n64) );
  INVX2 U68 ( .A(n108), .Y(n560) );
  INVX1 U69 ( .A(n552), .Y(n43) );
  OR2X2 U70 ( .A(n727), .B(n728), .Y(n504) );
  INVX1 U71 ( .A(n767), .Y(n79) );
  OR2X2 U72 ( .A(n722), .B(n82), .Y(n51) );
  AND2X2 U73 ( .A(\In<2> ), .B(n100), .Y(n44) );
  NOR2X1 U74 ( .A(n44), .B(n30), .Y(n638) );
  INVX1 U75 ( .A(n560), .Y(n45) );
  INVX1 U76 ( .A(n138), .Y(n92) );
  INVX2 U77 ( .A(n150), .Y(n62) );
  INVX1 U78 ( .A(n189), .Y(n47) );
  INVX1 U79 ( .A(n145), .Y(n48) );
  INVX1 U80 ( .A(n116), .Y(n117) );
  INVX1 U81 ( .A(n606), .Y(n49) );
  INVX1 U82 ( .A(\Cnt<1> ), .Y(n50) );
  OR2X2 U83 ( .A(n559), .B(n136), .Y(n353) );
  INVX1 U84 ( .A(n147), .Y(n102) );
  INVX1 U85 ( .A(n191), .Y(n578) );
  INVX1 U86 ( .A(n51), .Y(n52) );
  OR2X2 U87 ( .A(n86), .B(n87), .Y(n53) );
  INVX1 U88 ( .A(n53), .Y(n54) );
  OR2X2 U89 ( .A(n91), .B(n742), .Y(n55) );
  INVX1 U90 ( .A(n55), .Y(n56) );
  INVX1 U91 ( .A(n57), .Y(n58) );
  AND2X2 U92 ( .A(n526), .B(n319), .Y(n59) );
  AND2X2 U93 ( .A(n38), .B(n144), .Y(n426) );
  INVX1 U94 ( .A(n166), .Y(n60) );
  AND2X2 U95 ( .A(n29), .B(n574), .Y(n411) );
  AND2X2 U96 ( .A(n740), .B(n763), .Y(n561) );
  AND2X2 U97 ( .A(\In<9> ), .B(n139), .Y(n61) );
  INVX1 U98 ( .A(n61), .Y(n88) );
  OR2X2 U99 ( .A(n706), .B(n705), .Y(n501) );
  INVX2 U100 ( .A(n589), .Y(n590) );
  INVX4 U101 ( .A(n624), .Y(n768) );
  INVX1 U102 ( .A(n602), .Y(n95) );
  INVX1 U103 ( .A(n768), .Y(n78) );
  INVX1 U104 ( .A(n150), .Y(n151) );
  INVX1 U105 ( .A(n622), .Y(n614) );
  INVX1 U106 ( .A(n598), .Y(n65) );
  INVX1 U107 ( .A(n598), .Y(n749) );
  INVX1 U108 ( .A(n591), .Y(n606) );
  INVX1 U109 ( .A(n288), .Y(n67) );
  INVX1 U110 ( .A(\In<12> ), .Y(n69) );
  INVX1 U111 ( .A(n69), .Y(n70) );
  INVX1 U112 ( .A(n348), .Y(n71) );
  INVX1 U113 ( .A(n138), .Y(n72) );
  INVX1 U114 ( .A(n268), .Y(n589) );
  OR2X2 U115 ( .A(n717), .B(n718), .Y(n363) );
  OAI21X1 U116 ( .A(n62), .B(n269), .C(n468), .Y(n73) );
  INVX1 U117 ( .A(n397), .Y(n74) );
  INVX1 U118 ( .A(n160), .Y(n701) );
  BUFX2 U119 ( .A(n751), .Y(n75) );
  INVX1 U120 ( .A(n186), .Y(n76) );
  OR2X2 U121 ( .A(n761), .B(n760), .Y(n381) );
  INVX1 U122 ( .A(n167), .Y(n595) );
  OAI21X1 U123 ( .A(n78), .B(n79), .C(n464), .Y(n77) );
  INVX1 U124 ( .A(n77), .Y(n769) );
  INVX1 U125 ( .A(n615), .Y(n80) );
  NOR3X1 U126 ( .A(n73), .B(n469), .C(n363), .Y(n81) );
  INVX2 U127 ( .A(n120), .Y(n321) );
  OR2X1 U128 ( .A(n666), .B(n667), .Y(n246) );
  AND2X2 U129 ( .A(n763), .B(n751), .Y(n82) );
  INVX1 U130 ( .A(\In<9> ), .Y(n661) );
  BUFX4 U131 ( .A(n527), .Y(n588) );
  OR2X2 U132 ( .A(n137), .B(\Op<1> ), .Y(n83) );
  INVX1 U133 ( .A(n599), .Y(n84) );
  INVX1 U134 ( .A(n168), .Y(n85) );
  INVX2 U135 ( .A(n137), .Y(n764) );
  AND2X2 U136 ( .A(n104), .B(\In<10> ), .Y(n86) );
  AND2X2 U137 ( .A(\In<11> ), .B(n611), .Y(n87) );
  INVX1 U138 ( .A(n564), .Y(n109) );
  INVX1 U139 ( .A(\Cnt<1> ), .Y(n89) );
  NOR3X1 U140 ( .A(n320), .B(n174), .C(n264), .Y(n90) );
  AND2X2 U141 ( .A(n744), .B(n743), .Y(n91) );
  INVX1 U142 ( .A(n138), .Y(n139) );
  INVX1 U143 ( .A(n192), .Y(n93) );
  INVX1 U144 ( .A(\In<0> ), .Y(n671) );
  INVX8 U145 ( .A(n353), .Y(n757) );
  INVX1 U146 ( .A(n580), .Y(n579) );
  OAI21X1 U147 ( .A(n136), .B(n576), .C(n90), .Y(n94) );
  INVX1 U148 ( .A(n94), .Y(n660) );
  AND2X2 U149 ( .A(n144), .B(n588), .Y(n377) );
  AND2X2 U150 ( .A(n560), .B(n144), .Y(n421) );
  AND2X2 U151 ( .A(n144), .B(n190), .Y(n496) );
  INVX2 U152 ( .A(n645), .Y(n700) );
  INVX1 U153 ( .A(n622), .Y(n613) );
  OR2X2 U154 ( .A(n151), .B(n559), .Y(n143) );
  INVX1 U155 ( .A(\In<15> ), .Y(n657) );
  AND2X2 U156 ( .A(n46), .B(n753), .Y(n366) );
  AND2X2 U157 ( .A(n572), .B(n763), .Y(n391) );
  AND2X2 U158 ( .A(n764), .B(n33), .Y(n298) );
  AND2X2 U159 ( .A(n557), .B(n764), .Y(n545) );
  MUX2X1 U160 ( .B(n564), .A(n155), .S(n95), .Y(n744) );
  AND2X2 U161 ( .A(n726), .B(n37), .Y(n407) );
  OR2X2 U162 ( .A(n703), .B(n702), .Y(n356) );
  OR2X2 U163 ( .A(n83), .B(n192), .Y(n466) );
  OR2X2 U164 ( .A(n155), .B(n83), .Y(n468) );
  AND2X2 U165 ( .A(n24), .B(n741), .Y(n345) );
  INVX1 U166 ( .A(n187), .Y(n96) );
  OAI21X1 U167 ( .A(n41), .B(n661), .C(n7), .Y(n97) );
  INVX1 U168 ( .A(n97), .Y(n686) );
  INVX1 U169 ( .A(n164), .Y(n98) );
  AND2X2 U170 ( .A(n744), .B(n455), .Y(n355) );
  INVX1 U171 ( .A(\Cnt<2> ), .Y(n99) );
  INVX8 U172 ( .A(n321), .Y(n739) );
  INVX1 U173 ( .A(n147), .Y(n100) );
  INVX1 U174 ( .A(n147), .Y(n101) );
  INVX1 U175 ( .A(n147), .Y(n103) );
  INVX1 U176 ( .A(n147), .Y(n104) );
  INVX1 U177 ( .A(n102), .Y(n105) );
  INVX1 U178 ( .A(n520), .Y(n106) );
  AND2X2 U179 ( .A(\In<2> ), .B(n36), .Y(n294) );
  AND2X2 U180 ( .A(n560), .B(n753), .Y(n107) );
  AND2X2 U181 ( .A(n726), .B(n567), .Y(n420) );
  AND2X2 U182 ( .A(n757), .B(n566), .Y(n369) );
  NOR3X1 U183 ( .A(n525), .B(n109), .C(n499), .Y(n108) );
  NOR3X1 U184 ( .A(n61), .B(n354), .C(n551), .Y(n110) );
  AND2X2 U185 ( .A(n584), .B(n567), .Y(n403) );
  INVX1 U186 ( .A(n398), .Y(n114) );
  INVX1 U187 ( .A(n140), .Y(n111) );
  AND2X2 U188 ( .A(n111), .B(n267), .Y(n373) );
  AND2X2 U189 ( .A(n569), .B(n757), .Y(n413) );
  AND2X2 U190 ( .A(n569), .B(n753), .Y(n375) );
  INVX1 U191 ( .A(n158), .Y(n112) );
  NOR3X1 U192 ( .A(n114), .B(n272), .C(n4), .Y(n113) );
  AND2X2 U193 ( .A(n459), .B(n63), .Y(n378) );
  AND2X2 U194 ( .A(n768), .B(n572), .Y(n393) );
  AND2X2 U195 ( .A(n515), .B(n157), .Y(n634) );
  INVX1 U196 ( .A(n139), .Y(n682) );
  AND2X2 U197 ( .A(\In<15> ), .B(n80), .Y(n284) );
  AND2X2 U198 ( .A(n511), .B(n533), .Y(n659) );
  AND2X2 U199 ( .A(\In<14> ), .B(n607), .Y(n520) );
  AND2X2 U200 ( .A(n763), .B(n12), .Y(n494) );
  AND2X2 U201 ( .A(n451), .B(n352), .Y(n115) );
  AND2X2 U202 ( .A(n535), .B(n134), .Y(n116) );
  OR2X2 U203 ( .A(n606), .B(n601), .Y(n118) );
  OR2X2 U204 ( .A(n670), .B(n136), .Y(n119) );
  INVX1 U205 ( .A(n119), .Y(n120) );
  OR2X2 U206 ( .A(n632), .B(n137), .Y(n121) );
  OR2X2 U207 ( .A(n632), .B(n151), .Y(n122) );
  INVX1 U208 ( .A(n122), .Y(n123) );
  AND2X2 U209 ( .A(n660), .B(n245), .Y(n124) );
  INVX1 U210 ( .A(n124), .Y(\Out<1> ) );
  AND2X2 U211 ( .A(n247), .B(n678), .Y(n126) );
  INVX1 U212 ( .A(n126), .Y(\Out<2> ) );
  OR2X2 U213 ( .A(n462), .B(n711), .Y(n128) );
  INVX1 U214 ( .A(n128), .Y(n129) );
  AND2X2 U215 ( .A(\In<4> ), .B(n103), .Y(n130) );
  OR2X2 U216 ( .A(n522), .B(n351), .Y(\Out<4> ) );
  AND2X2 U217 ( .A(n133), .B(n304), .Y(n132) );
  AND2X2 U218 ( .A(n542), .B(n5), .Y(n133) );
  AND2X2 U219 ( .A(n524), .B(n347), .Y(n134) );
  OR2X2 U220 ( .A(n624), .B(n586), .Y(n135) );
  OR2X2 U221 ( .A(n66), .B(n600), .Y(n136) );
  OR2X2 U222 ( .A(n66), .B(\Cnt<3> ), .Y(n137) );
  OR2X2 U223 ( .A(\Cnt<1> ), .B(\Cnt<0> ), .Y(n138) );
  AND2X2 U224 ( .A(n596), .B(n597), .Y(n140) );
  OR2X2 U225 ( .A(n25), .B(n599), .Y(n141) );
  INVX1 U226 ( .A(n141), .Y(n142) );
  INVX1 U227 ( .A(n143), .Y(n144) );
  AND2X2 U228 ( .A(n656), .B(n655), .Y(n145) );
  INVX1 U229 ( .A(n145), .Y(n146) );
  OR2X2 U230 ( .A(n89), .B(\Cnt<0> ), .Y(n147) );
  INVX1 U231 ( .A(n147), .Y(n148) );
  OR2X2 U232 ( .A(n62), .B(n670), .Y(n149) );
  AND2X2 U233 ( .A(\Cnt<3> ), .B(n99), .Y(n150) );
  AND2X2 U234 ( .A(n54), .B(n237), .Y(n152) );
  AND2X2 U235 ( .A(n300), .B(n439), .Y(n153) );
  INVX1 U236 ( .A(n153), .Y(n154) );
  AND2X2 U237 ( .A(n302), .B(n441), .Y(n155) );
  AND2X2 U238 ( .A(\In<15> ), .B(n612), .Y(n156) );
  INVX1 U239 ( .A(n156), .Y(n157) );
  AND2X2 U240 ( .A(n634), .B(n238), .Y(n158) );
  AND2X2 U241 ( .A(n715), .B(n764), .Y(n159) );
  INVX1 U242 ( .A(n159), .Y(n160) );
  AND2X2 U243 ( .A(\In<11> ), .B(n616), .Y(n161) );
  AND2X2 U244 ( .A(n449), .B(n432), .Y(n162) );
  AND2X2 U245 ( .A(\In<3> ), .B(n612), .Y(n163) );
  AND2X2 U246 ( .A(n434), .B(n312), .Y(n164) );
  AND2X2 U247 ( .A(n103), .B(\In<11> ), .Y(n324) );
  AND2X2 U248 ( .A(\In<10> ), .B(n607), .Y(n165) );
  AND2X2 U249 ( .A(n148), .B(\In<7> ), .Y(n166) );
  OR2X2 U250 ( .A(n261), .B(n249), .Y(n167) );
  AND2X2 U251 ( .A(\In<5> ), .B(n68), .Y(n168) );
  AND2X2 U252 ( .A(n648), .B(n647), .Y(n169) );
  AND2X2 U253 ( .A(n653), .B(n654), .Y(n170) );
  AND2X2 U254 ( .A(\In<4> ), .B(n609), .Y(n171) );
  INVX1 U255 ( .A(n171), .Y(n172) );
  AND2X2 U256 ( .A(\In<1> ), .B(n92), .Y(n173) );
  AND2X2 U257 ( .A(n726), .B(n146), .Y(n174) );
  AND2X2 U258 ( .A(\In<10> ), .B(n92), .Y(n176) );
  AND2X2 U259 ( .A(\In<12> ), .B(n101), .Y(n177) );
  AND2X2 U260 ( .A(n664), .B(n239), .Y(n178) );
  AND2X2 U261 ( .A(n557), .B(n669), .Y(n179) );
  INVX1 U262 ( .A(n179), .Y(n180) );
  AND2X2 U263 ( .A(n242), .B(n180), .Y(n181) );
  OR2X2 U264 ( .A(n157), .B(n670), .Y(n182) );
  AND2X2 U265 ( .A(n675), .B(n674), .Y(n183) );
  INVX1 U266 ( .A(n183), .Y(n184) );
  AND2X2 U267 ( .A(n443), .B(n306), .Y(n185) );
  AND2X2 U268 ( .A(n683), .B(n281), .Y(n186) );
  AND2X2 U269 ( .A(n686), .B(n436), .Y(n187) );
  INVX1 U270 ( .A(n187), .Y(n188) );
  AND2X2 U271 ( .A(n314), .B(n240), .Y(n189) );
  INVX1 U272 ( .A(n189), .Y(n190) );
  AND2X2 U273 ( .A(n308), .B(n445), .Y(n191) );
  AND2X2 U274 ( .A(n243), .B(n310), .Y(n192) );
  INVX1 U275 ( .A(n192), .Y(n193) );
  AND2X2 U276 ( .A(n584), .B(n570), .Y(n194) );
  INVX1 U277 ( .A(n194), .Y(n195) );
  AND2X2 U278 ( .A(n184), .B(n741), .Y(n196) );
  OR2X2 U279 ( .A(n317), .B(n342), .Y(n197) );
  AND2X2 U280 ( .A(n768), .B(n539), .Y(n198) );
  INVX1 U281 ( .A(n198), .Y(n199) );
  AND2X2 U282 ( .A(n587), .B(n651), .Y(n200) );
  INVX1 U283 ( .A(n200), .Y(n201) );
  AND2X2 U284 ( .A(n762), .B(n571), .Y(n202) );
  INVX1 U285 ( .A(n202), .Y(n203) );
  AND2X2 U286 ( .A(n585), .B(n350), .Y(n204) );
  INVX1 U287 ( .A(n204), .Y(n205) );
  INVX1 U288 ( .A(n209), .Y(n206) );
  AND2X2 U289 ( .A(n123), .B(n14), .Y(n207) );
  INVX1 U290 ( .A(n207), .Y(n208) );
  AND2X2 U291 ( .A(n100), .B(\In<8> ), .Y(n209) );
  AND2X2 U292 ( .A(n523), .B(n71), .Y(n210) );
  INVX1 U293 ( .A(n210), .Y(n211) );
  AND2X2 U294 ( .A(n740), .B(n672), .Y(n212) );
  AND2X2 U295 ( .A(n144), .B(n76), .Y(n213) );
  INVX1 U296 ( .A(n213), .Y(n214) );
  AND2X2 U297 ( .A(n739), .B(n536), .Y(n215) );
  INVX1 U298 ( .A(n215), .Y(n216) );
  AND2X2 U299 ( .A(n585), .B(n577), .Y(n217) );
  INVX1 U300 ( .A(n217), .Y(n218) );
  AND2X2 U301 ( .A(n701), .B(n111), .Y(n219) );
  INVX1 U302 ( .A(n219), .Y(n220) );
  AND2X2 U303 ( .A(n584), .B(n38), .Y(n221) );
  INVX1 U304 ( .A(n221), .Y(n222) );
  AND2X2 U305 ( .A(n584), .B(n527), .Y(n223) );
  INVX1 U306 ( .A(n223), .Y(n224) );
  AND2X2 U307 ( .A(n701), .B(n573), .Y(n225) );
  INVX1 U308 ( .A(n225), .Y(n226) );
  AND2X2 U309 ( .A(\In<0> ), .B(n148), .Y(n227) );
  INVX1 U310 ( .A(n227), .Y(n228) );
  AND2X2 U311 ( .A(n726), .B(n568), .Y(n229) );
  INVX1 U312 ( .A(n229), .Y(n230) );
  AND2X2 U313 ( .A(n584), .B(n188), .Y(n231) );
  INVX1 U314 ( .A(n231), .Y(n232) );
  AND2X2 U315 ( .A(n739), .B(n24), .Y(n233) );
  INVX1 U316 ( .A(n233), .Y(n234) );
  AND2X2 U317 ( .A(n267), .B(n93), .Y(n235) );
  INVX1 U318 ( .A(n235), .Y(n236) );
  BUFX2 U319 ( .A(n626), .Y(n237) );
  BUFX2 U320 ( .A(n633), .Y(n238) );
  BUFX2 U321 ( .A(n665), .Y(n239) );
  BUFX2 U322 ( .A(n689), .Y(n240) );
  AND2X2 U323 ( .A(n587), .B(n211), .Y(n241) );
  INVX1 U324 ( .A(n241), .Y(n242) );
  BUFX2 U325 ( .A(n695), .Y(n243) );
  OR2X2 U326 ( .A(n650), .B(n649), .Y(n244) );
  INVX1 U327 ( .A(n244), .Y(n245) );
  INVX1 U328 ( .A(n246), .Y(n247) );
  AND2X2 U329 ( .A(n60), .B(n118), .Y(n248) );
  INVX1 U330 ( .A(n248), .Y(n249) );
  AND2X2 U331 ( .A(n199), .B(n208), .Y(n250) );
  INVX1 U332 ( .A(n250), .Y(n251) );
  AND2X2 U333 ( .A(n206), .B(n453), .Y(n252) );
  INVX1 U334 ( .A(n252), .Y(n253) );
  AND2X2 U335 ( .A(n543), .B(n517), .Y(n254) );
  INVX1 U336 ( .A(n254), .Y(n255) );
  INVX1 U337 ( .A(n256), .Y(n257) );
  AND2X2 U338 ( .A(n513), .B(n206), .Y(n258) );
  INVX1 U339 ( .A(n258), .Y(n259) );
  AND2X2 U340 ( .A(n141), .B(n88), .Y(n260) );
  INVX1 U341 ( .A(n260), .Y(n261) );
  OR2X2 U342 ( .A(n251), .B(n631), .Y(n262) );
  INVX1 U343 ( .A(n262), .Y(n263) );
  AND2X2 U344 ( .A(n553), .B(n739), .Y(n264) );
  OR2X2 U345 ( .A(n257), .B(n687), .Y(n265) );
  INVX1 U346 ( .A(n265), .Y(n266) );
  AND2X2 U347 ( .A(n740), .B(n768), .Y(n267) );
  INVX1 U348 ( .A(n267), .Y(n268) );
  AND2X2 U349 ( .A(n540), .B(n362), .Y(n269) );
  BUFX2 U350 ( .A(n644), .Y(n270) );
  BUFX2 U351 ( .A(n698), .Y(n271) );
  AND2X2 U352 ( .A(n101), .B(\In<15> ), .Y(n272) );
  BUFX2 U353 ( .A(n643), .Y(n273) );
  OR2X2 U354 ( .A(n696), .B(n697), .Y(n274) );
  INVX1 U355 ( .A(n274), .Y(n275) );
  AND2X2 U356 ( .A(\In<3> ), .B(n102), .Y(n276) );
  INVX1 U357 ( .A(n276), .Y(n277) );
  INVX1 U358 ( .A(n276), .Y(n278) );
  AND2X2 U359 ( .A(\In<13> ), .B(n148), .Y(n279) );
  INVX1 U360 ( .A(n279), .Y(n280) );
  AND2X2 U361 ( .A(n521), .B(n280), .Y(n281) );
  INVX1 U362 ( .A(n281), .Y(n282) );
  AND2X2 U363 ( .A(\In<14> ), .B(n104), .Y(n283) );
  AND2X2 U364 ( .A(\In<7> ), .B(n18), .Y(n285) );
  AND2X2 U365 ( .A(n616), .B(\In<6> ), .Y(n286) );
  INVX1 U366 ( .A(n286), .Y(n287) );
  AND2X2 U367 ( .A(\In<2> ), .B(n611), .Y(n288) );
  AND2X2 U368 ( .A(\In<4> ), .B(n617), .Y(n289) );
  AND2X2 U369 ( .A(\In<6> ), .B(n139), .Y(n290) );
  AND2X2 U370 ( .A(\In<12> ), .B(n618), .Y(n291) );
  INVX1 U371 ( .A(n291), .Y(n292) );
  INVX1 U372 ( .A(n197), .Y(n293) );
  INVX1 U373 ( .A(n294), .Y(n295) );
  AND2X2 U374 ( .A(\In<5> ), .B(n617), .Y(n296) );
  INVX1 U375 ( .A(n296), .Y(n297) );
  INVX1 U376 ( .A(n298), .Y(n299) );
  BUFX2 U377 ( .A(n627), .Y(n300) );
  INVX1 U378 ( .A(n629), .Y(n301) );
  INVX1 U379 ( .A(n301), .Y(n302) );
  INVX1 U380 ( .A(n676), .Y(n303) );
  INVX1 U381 ( .A(n303), .Y(n304) );
  INVX1 U382 ( .A(n679), .Y(n305) );
  INVX1 U383 ( .A(n305), .Y(n306) );
  INVX1 U384 ( .A(n691), .Y(n307) );
  INVX1 U385 ( .A(n307), .Y(n308) );
  INVX1 U386 ( .A(n694), .Y(n309) );
  INVX1 U387 ( .A(n309), .Y(n310) );
  INVX1 U388 ( .A(n640), .Y(n311) );
  INVX1 U389 ( .A(n311), .Y(n312) );
  INVX1 U390 ( .A(n690), .Y(n313) );
  INVX1 U391 ( .A(n313), .Y(n314) );
  INVX1 U392 ( .A(n110), .Y(n315) );
  INVX1 U393 ( .A(n733), .Y(n316) );
  INVX1 U394 ( .A(n316), .Y(n317) );
  INVX1 U395 ( .A(n684), .Y(n318) );
  INVX1 U396 ( .A(n318), .Y(n319) );
  AND2X2 U397 ( .A(n768), .B(n751), .Y(n320) );
  INVX1 U398 ( .A(n120), .Y(n322) );
  INVX1 U399 ( .A(n105), .Y(n323) );
  INVX1 U400 ( .A(\In<6> ), .Y(n601) );
  AND2X2 U401 ( .A(n757), .B(n338), .Y(n325) );
  INVX1 U402 ( .A(n325), .Y(n326) );
  AND2X2 U403 ( .A(n741), .B(n6), .Y(n327) );
  AND2X2 U404 ( .A(n757), .B(n570), .Y(n328) );
  INVX1 U405 ( .A(n328), .Y(n329) );
  INVX1 U406 ( .A(n324), .Y(n330) );
  AND2X2 U407 ( .A(\In<8> ), .B(n610), .Y(n331) );
  INVX1 U408 ( .A(n331), .Y(n332) );
  INVX1 U409 ( .A(n334), .Y(n333) );
  INVX1 U410 ( .A(n327), .Y(n335) );
  INVX1 U411 ( .A(n196), .Y(n336) );
  INVX1 U412 ( .A(n166), .Y(n337) );
  INVX1 U413 ( .A(n145), .Y(n338) );
  INVX1 U414 ( .A(n772), .Y(n339) );
  INVX1 U415 ( .A(n339), .Y(\Out<13> ) );
  INVX1 U416 ( .A(n734), .Y(n341) );
  INVX1 U417 ( .A(n341), .Y(n342) );
  INVX1 U418 ( .A(n343), .Y(n344) );
  INVX1 U419 ( .A(n345), .Y(n346) );
  INVX1 U420 ( .A(n283), .Y(n347) );
  AND2X2 U421 ( .A(n139), .B(\In<14> ), .Y(n348) );
  INVX1 U422 ( .A(n348), .Y(n349) );
  INVX1 U423 ( .A(n185), .Y(n350) );
  INVX1 U424 ( .A(n587), .Y(n632) );
  OR2X2 U425 ( .A(n356), .B(n355), .Y(n351) );
  INVX1 U426 ( .A(\In<8> ), .Y(n599) );
  AND2X2 U427 ( .A(\In<10> ), .B(n619), .Y(n354) );
  AND2X2 U428 ( .A(n457), .B(n195), .Y(n357) );
  INVX1 U429 ( .A(n357), .Y(n358) );
  AND2X2 U430 ( .A(n726), .B(n96), .Y(n359) );
  INVX1 U431 ( .A(n359), .Y(n360) );
  AND2X2 U432 ( .A(n715), .B(n117), .Y(n361) );
  INVX1 U433 ( .A(n361), .Y(n362) );
  AND2X2 U434 ( .A(n739), .B(n565), .Y(n364) );
  AND2X2 U435 ( .A(n144), .B(n569), .Y(n365) );
  AND2X2 U436 ( .A(n98), .B(n741), .Y(n367) );
  INVX1 U437 ( .A(n367), .Y(n368) );
  AND2X2 U438 ( .A(n48), .B(n753), .Y(n370) );
  INVX1 U439 ( .A(n370), .Y(n371) );
  INVX1 U440 ( .A(n373), .Y(n374) );
  INVX1 U441 ( .A(n375), .Y(n376) );
  INVX1 U442 ( .A(n546), .Y(n753) );
  AND2X2 U443 ( .A(n144), .B(n96), .Y(n379) );
  INVX1 U444 ( .A(n379), .Y(n380) );
  INVX1 U445 ( .A(n381), .Y(n382) );
  INVX1 U446 ( .A(n652), .Y(n383) );
  INVX1 U447 ( .A(n383), .Y(n384) );
  INVX1 U448 ( .A(n21), .Y(\Out<5> ) );
  INVX1 U449 ( .A(n279), .Y(n387) );
  INVX1 U450 ( .A(n161), .Y(n388) );
  OR2X1 U451 ( .A(n710), .B(n709), .Y(n389) );
  INVX1 U452 ( .A(n389), .Y(n390) );
  INVX1 U453 ( .A(n391), .Y(n392) );
  INVX1 U454 ( .A(n393), .Y(n394) );
  AND2X2 U455 ( .A(n382), .B(n769), .Y(n395) );
  INVX1 U456 ( .A(n395), .Y(\Out<15> ) );
  AND2X2 U457 ( .A(n18), .B(\In<14> ), .Y(n397) );
  INVX1 U458 ( .A(n397), .Y(n398) );
  INVX1 U459 ( .A(n291), .Y(n399) );
  INVX1 U460 ( .A(n175), .Y(n400) );
  AND2X2 U461 ( .A(\In<2> ), .B(n72), .Y(n401) );
  INVX1 U462 ( .A(n401), .Y(n402) );
  INVX1 U463 ( .A(n403), .Y(n404) );
  AND2X2 U464 ( .A(n554), .B(n585), .Y(n405) );
  INVX1 U465 ( .A(n405), .Y(n406) );
  INVX1 U466 ( .A(n407), .Y(n408) );
  AND2X2 U467 ( .A(n585), .B(n111), .Y(n409) );
  INVX1 U468 ( .A(n409), .Y(n410) );
  INVX1 U469 ( .A(n411), .Y(n412) );
  INVX1 U470 ( .A(n413), .Y(n414) );
  AND2X1 U471 ( .A(n726), .B(n588), .Y(n415) );
  INVX1 U472 ( .A(n415), .Y(n416) );
  AND2X1 U473 ( .A(n736), .B(n580), .Y(n417) );
  INVX1 U474 ( .A(n417), .Y(n418) );
  INVX1 U475 ( .A(n420), .Y(n419) );
  INVX1 U476 ( .A(n421), .Y(n422) );
  INVX1 U477 ( .A(n364), .Y(n423) );
  INVX1 U478 ( .A(n365), .Y(n424) );
  INVX1 U479 ( .A(n369), .Y(n425) );
  INVX1 U480 ( .A(n426), .Y(n427) );
  AND2X1 U481 ( .A(n574), .B(n267), .Y(n428) );
  INVX1 U482 ( .A(n428), .Y(n429) );
  INVX1 U483 ( .A(n377), .Y(n430) );
  INVX1 U484 ( .A(n636), .Y(n431) );
  INVX1 U485 ( .A(n431), .Y(n432) );
  INVX1 U486 ( .A(n639), .Y(n433) );
  INVX1 U487 ( .A(n433), .Y(n434) );
  INVX1 U488 ( .A(n685), .Y(n435) );
  INVX1 U489 ( .A(n435), .Y(n436) );
  INVX1 U490 ( .A(n130), .Y(n437) );
  INVX1 U491 ( .A(n628), .Y(n438) );
  INVX1 U492 ( .A(n438), .Y(n439) );
  INVX1 U493 ( .A(n630), .Y(n440) );
  INVX1 U494 ( .A(n440), .Y(n441) );
  INVX1 U495 ( .A(n680), .Y(n442) );
  INVX1 U496 ( .A(n442), .Y(n443) );
  INVX1 U497 ( .A(n692), .Y(n444) );
  INVX1 U498 ( .A(n444), .Y(n445) );
  INVX1 U499 ( .A(n738), .Y(n446) );
  INVX1 U500 ( .A(n446), .Y(n447) );
  INVX1 U501 ( .A(n637), .Y(n448) );
  INVX1 U502 ( .A(n448), .Y(n449) );
  INVX1 U503 ( .A(n737), .Y(n450) );
  INVX1 U504 ( .A(n450), .Y(n451) );
  AND2X2 U505 ( .A(\In<7> ), .B(n607), .Y(n452) );
  INVX1 U506 ( .A(n452), .Y(n453) );
  OR2X1 U507 ( .A(n603), .B(\Op<1> ), .Y(n454) );
  INVX1 U508 ( .A(n454), .Y(n455) );
  AND2X2 U509 ( .A(n739), .B(n10), .Y(n456) );
  INVX1 U510 ( .A(n456), .Y(n457) );
  OR2X1 U511 ( .A(n755), .B(n754), .Y(n458) );
  INVX1 U512 ( .A(n458), .Y(n459) );
  INVX1 U513 ( .A(n378), .Y(\Out<14> ) );
  AND2X2 U514 ( .A(n392), .B(n299), .Y(n461) );
  INVX1 U515 ( .A(n461), .Y(n462) );
  AND2X2 U516 ( .A(n394), .B(n333), .Y(n463) );
  INVX1 U517 ( .A(n766), .Y(n464) );
  INVX1 U518 ( .A(n182), .Y(n465) );
  INVX1 U519 ( .A(n466), .Y(n467) );
  INVX1 U520 ( .A(n470), .Y(n469) );
  BUFX2 U521 ( .A(n719), .Y(n470) );
  BUFX2 U522 ( .A(n730), .Y(n471) );
  BUFX2 U523 ( .A(n746), .Y(n472) );
  INVX1 U524 ( .A(n474), .Y(n473) );
  BUFX2 U525 ( .A(n708), .Y(n474) );
  INVX1 U526 ( .A(n714), .Y(n475) );
  INVX1 U527 ( .A(n475), .Y(n476) );
  BUFX2 U528 ( .A(n724), .Y(n477) );
  AND2X2 U529 ( .A(n267), .B(n10), .Y(n478) );
  INVX1 U530 ( .A(n478), .Y(n479) );
  AND2X2 U531 ( .A(n764), .B(n350), .Y(n480) );
  INVX1 U532 ( .A(n480), .Y(n481) );
  INVX1 U533 ( .A(n765), .Y(n482) );
  INVX1 U534 ( .A(n482), .Y(n483) );
  BUFX2 U535 ( .A(n773), .Y(\Out<7> ) );
  INVX1 U536 ( .A(n486), .Y(\Out<6> ) );
  AND2X2 U537 ( .A(n390), .B(n129), .Y(n486) );
  OR2X2 U538 ( .A(n282), .B(n688), .Y(n487) );
  INVX1 U539 ( .A(n487), .Y(n488) );
  OR2X1 U540 ( .A(n136), .B(n632), .Y(n489) );
  INVX1 U541 ( .A(n489), .Y(n490) );
  BUFX2 U542 ( .A(n713), .Y(n491) );
  BUFX2 U543 ( .A(n729), .Y(n492) );
  BUFX2 U544 ( .A(n723), .Y(n493) );
  INVX1 U545 ( .A(n496), .Y(n495) );
  AND2X2 U546 ( .A(n768), .B(n12), .Y(n497) );
  INVX1 U547 ( .A(n497), .Y(n498) );
  INVX1 U548 ( .A(n638), .Y(n499) );
  BUFX2 U549 ( .A(n752), .Y(n500) );
  OR2X2 U550 ( .A(n358), .B(n712), .Y(n502) );
  INVX1 U551 ( .A(n502), .Y(n503) );
  INVX1 U552 ( .A(n504), .Y(n505) );
  INVX1 U553 ( .A(n366), .Y(n506) );
  AND2X2 U554 ( .A(n757), .B(n96), .Y(n507) );
  INVX1 U555 ( .A(n507), .Y(n508) );
  INVX1 U556 ( .A(n165), .Y(n509) );
  INVX1 U557 ( .A(n168), .Y(n510) );
  INVX1 U558 ( .A(n173), .Y(n511) );
  AND2X2 U559 ( .A(\In<9> ), .B(n609), .Y(n512) );
  INVX1 U560 ( .A(n512), .Y(n513) );
  INVX1 U561 ( .A(n512), .Y(n514) );
  INVX1 U562 ( .A(n283), .Y(n515) );
  INVX1 U563 ( .A(n290), .Y(n516) );
  INVX1 U564 ( .A(n290), .Y(n517) );
  INVX1 U565 ( .A(n176), .Y(n518) );
  INVX1 U566 ( .A(n118), .Y(n519) );
  INVX1 U567 ( .A(n520), .Y(n521) );
  INVX1 U568 ( .A(n704), .Y(n522) );
  INVX1 U569 ( .A(n284), .Y(n523) );
  INVX1 U570 ( .A(n284), .Y(n524) );
  INVX1 U571 ( .A(n28), .Y(n525) );
  INVX1 U572 ( .A(n288), .Y(n526) );
  OR2X2 U573 ( .A(n259), .B(n255), .Y(n527) );
  INVX1 U574 ( .A(n527), .Y(n528) );
  AND2X2 U575 ( .A(n619), .B(\In<13> ), .Y(n529) );
  INVX1 U576 ( .A(n529), .Y(n530) );
  INVX1 U577 ( .A(n289), .Y(n531) );
  AND2X2 U578 ( .A(\In<0> ), .B(n36), .Y(n532) );
  INVX1 U579 ( .A(n9), .Y(n533) );
  AND2X2 U580 ( .A(\In<13> ), .B(n609), .Y(n534) );
  INVX1 U581 ( .A(n534), .Y(n535) );
  INVX1 U582 ( .A(n155), .Y(n536) );
  AND2X2 U583 ( .A(n92), .B(\In<13> ), .Y(n537) );
  INVX1 U584 ( .A(n537), .Y(n538) );
  AND2X2 U585 ( .A(n740), .B(n563), .Y(n539) );
  INVX1 U586 ( .A(n539), .Y(n540) );
  AND2X2 U587 ( .A(\In<5> ), .B(n612), .Y(n541) );
  INVX1 U588 ( .A(n541), .Y(n542) );
  INVX1 U589 ( .A(n285), .Y(n543) );
  INVX1 U590 ( .A(n115), .Y(\Out<11> ) );
  INVX1 U591 ( .A(n545), .Y(n546) );
  INVX1 U592 ( .A(n725), .Y(n547) );
  INVX1 U593 ( .A(n547), .Y(n548) );
  INVX1 U594 ( .A(n177), .Y(n549) );
  INVX1 U595 ( .A(n551), .Y(n550) );
  AND2X2 U596 ( .A(\In<12> ), .B(n608), .Y(n551) );
  INVX1 U597 ( .A(n758), .Y(n552) );
  INVX1 U598 ( .A(n731), .Y(n758) );
  INVX1 U599 ( .A(n170), .Y(n553) );
  INVX1 U600 ( .A(n162), .Y(n554) );
  AND2X2 U601 ( .A(\Op<1> ), .B(\Op<0> ), .Y(n555) );
  INVX1 U602 ( .A(n555), .Y(n556) );
  AND2X2 U603 ( .A(\Op<1> ), .B(n625), .Y(n557) );
  INVX1 U604 ( .A(n557), .Y(n558) );
  INVX1 U605 ( .A(n557), .Y(n559) );
  INVX1 U606 ( .A(n561), .Y(n562) );
  AND2X2 U607 ( .A(\In<0> ), .B(n68), .Y(n563) );
  INVX1 U608 ( .A(n563), .Y(n564) );
  INVX1 U609 ( .A(n140), .Y(n565) );
  INVX1 U610 ( .A(n152), .Y(n566) );
  INVX1 U611 ( .A(n152), .Y(n567) );
  INVX1 U612 ( .A(n132), .Y(n568) );
  INVX1 U613 ( .A(n132), .Y(n569) );
  INVX1 U614 ( .A(n1), .Y(n570) );
  INVX1 U615 ( .A(n181), .Y(n571) );
  INVX1 U616 ( .A(n181), .Y(n572) );
  INVX1 U617 ( .A(n178), .Y(n573) );
  INVX1 U618 ( .A(n178), .Y(n574) );
  INVX1 U619 ( .A(n576), .Y(n575) );
  AND2X2 U620 ( .A(n201), .B(n384), .Y(n576) );
  INVX1 U621 ( .A(n164), .Y(n577) );
  AND2X2 U622 ( .A(\In<15> ), .B(n68), .Y(n580) );
  INVX1 U623 ( .A(n580), .Y(n581) );
  OR2X2 U624 ( .A(n253), .B(n662), .Y(n583) );
  INVX1 U625 ( .A(\Op<0> ), .Y(n625) );
  AND2X2 U626 ( .A(n558), .B(n556), .Y(n586) );
  INVX1 U627 ( .A(n586), .Y(n587) );
  INVX2 U628 ( .A(n135), .Y(n726) );
  INVX1 U629 ( .A(n47), .Y(n759) );
  INVX1 U630 ( .A(n688), .Y(n683) );
  AND2X2 U631 ( .A(\Cnt<1> ), .B(\Cnt<0> ), .Y(n591) );
  OR2X2 U632 ( .A(n623), .B(n78), .Y(n592) );
  INVX1 U633 ( .A(n554), .Y(n716) );
  INVX1 U634 ( .A(n514), .Y(n635) );
  AND2X2 U635 ( .A(n592), .B(n593), .Y(n678) );
  AND2X2 U636 ( .A(n203), .B(n594), .Y(n593) );
  INVX1 U637 ( .A(n677), .Y(n594) );
  AND2X2 U638 ( .A(n509), .B(n330), .Y(n596) );
  AND2X2 U639 ( .A(n292), .B(n538), .Y(n597) );
  OR2X2 U640 ( .A(n315), .B(n646), .Y(n598) );
  INVX1 U641 ( .A(\In<11> ), .Y(n681) );
  INVX1 U642 ( .A(\Cnt<3> ), .Y(n600) );
  INVX1 U643 ( .A(n670), .Y(n715) );
  INVX1 U644 ( .A(n136), .Y(n762) );
  INVX1 U645 ( .A(n99), .Y(n602) );
  INVX1 U646 ( .A(n600), .Y(n603) );
  INVX1 U647 ( .A(n610), .Y(n604) );
  INVX1 U648 ( .A(n591), .Y(n605) );
  INVX1 U649 ( .A(n605), .Y(n607) );
  INVX1 U650 ( .A(n606), .Y(n608) );
  INVX1 U651 ( .A(n19), .Y(n609) );
  INVX1 U652 ( .A(n19), .Y(n610) );
  INVX1 U653 ( .A(n605), .Y(n611) );
  INVX1 U654 ( .A(n19), .Y(n612) );
  INVX1 U655 ( .A(n622), .Y(n615) );
  INVX1 U656 ( .A(n614), .Y(n616) );
  INVX1 U657 ( .A(n614), .Y(n617) );
  INVX1 U658 ( .A(n613), .Y(n618) );
  INVX1 U659 ( .A(n613), .Y(n619) );
  INVX1 U660 ( .A(n615), .Y(n620) );
  INVX1 U661 ( .A(n615), .Y(n621) );
  AND2X2 U662 ( .A(\Cnt<0> ), .B(n50), .Y(n622) );
  INVX1 U663 ( .A(n330), .Y(n646) );
  OR2X2 U664 ( .A(\Cnt<2> ), .B(\Cnt<3> ), .Y(n624) );
  INVX2 U665 ( .A(\Op<1> ), .Y(n740) );
  AOI22X1 U666 ( .A(n84), .B(n68), .C(\In<9> ), .D(n616), .Y(n626) );
  AOI22X1 U667 ( .A(\In<6> ), .B(n323), .C(\In<7> ), .D(n49), .Y(n628) );
  AOI22X1 U668 ( .A(\In<5> ), .B(n621), .C(\In<4> ), .D(n11), .Y(n627) );
  OR2X2 U669 ( .A(\Op<0> ), .B(\Op<1> ), .Y(n670) );
  AOI22X1 U670 ( .A(\In<2> ), .B(n23), .C(\In<1> ), .D(n608), .Y(n630) );
  AOI22X1 U671 ( .A(\In<3> ), .B(n620), .C(n20), .D(\In<4> ), .Y(n629) );
  OAI21X1 U672 ( .A(n153), .B(n121), .C(n216), .Y(n631) );
  AOI21X1 U673 ( .A(n70), .B(n72), .C(n529), .Y(n633) );
  AOI21X1 U674 ( .A(\In<10> ), .B(n31), .C(n635), .Y(n637) );
  AOI21X1 U675 ( .A(n70), .B(n72), .C(n161), .Y(n636) );
  AOI22X1 U676 ( .A(n490), .B(n112), .C(n701), .D(n27), .Y(n644) );
  AND2X2 U677 ( .A(n715), .B(n768), .Y(n642) );
  AOI21X1 U678 ( .A(\In<6> ), .B(n323), .C(n541), .Y(n640) );
  AOI21X1 U679 ( .A(\In<8> ), .B(n20), .C(n285), .Y(n639) );
  OAI21X1 U680 ( .A(n135), .B(n45), .C(n218), .Y(n641) );
  NAND3X1 U681 ( .A(n273), .B(n270), .C(n263), .Y(\Out<0> ) );
  OAI21X1 U682 ( .A(n556), .B(n151), .C(n143), .Y(n645) );
  OAI21X1 U683 ( .A(n749), .B(n700), .C(n220), .Y(n650) );
  AND2X2 U684 ( .A(n337), .B(n332), .Y(n648) );
  AND2X2 U685 ( .A(n85), .B(n287), .Y(n647) );
  OAI21X1 U686 ( .A(n22), .B(n149), .C(n222), .Y(n649) );
  NAND3X1 U687 ( .A(\In<0> ), .B(n557), .C(n608), .Y(n652) );
  AND2X2 U688 ( .A(n67), .B(n278), .Y(n654) );
  AND2X2 U689 ( .A(n531), .B(n510), .Y(n653) );
  AND2X2 U690 ( .A(n277), .B(n172), .Y(n656) );
  AND2X2 U691 ( .A(n511), .B(n295), .Y(n655) );
  OAI21X1 U692 ( .A(n13), .B(n657), .C(n106), .Y(n658) );
  OAI21X1 U693 ( .A(n659), .B(\Op<1> ), .C(n400), .Y(n751) );
  OAI21X1 U694 ( .A(n8), .B(n661), .C(n518), .Y(n662) );
  OAI21X1 U695 ( .A(n582), .B(n149), .C(n224), .Y(n667) );
  AND2X2 U696 ( .A(n388), .B(n518), .Y(n663) );
  NAND3X1 U697 ( .A(n535), .B(n549), .C(n663), .Y(n725) );
  AOI21X1 U698 ( .A(\In<11> ), .B(n49), .C(n177), .Y(n665) );
  AND2X2 U699 ( .A(n349), .B(n530), .Y(n664) );
  OAI21X1 U700 ( .A(n547), .B(n700), .C(n226), .Y(n666) );
  OAI21X1 U701 ( .A(n604), .B(n668), .C(n228), .Y(n669) );
  AOI21X1 U702 ( .A(n740), .B(n30), .C(n465), .Y(n673) );
  OAI21X1 U703 ( .A(n41), .B(n671), .C(n402), .Y(n672) );
  AND2X2 U704 ( .A(n437), .B(n28), .Y(n675) );
  AND2X2 U705 ( .A(n516), .B(n297), .Y(n674) );
  AOI22X1 U706 ( .A(\In<3> ), .B(n620), .C(\In<2> ), .D(n72), .Y(n676) );
  OAI21X1 U707 ( .A(n183), .B(n322), .C(n230), .Y(n677) );
  AOI22X1 U708 ( .A(\In<9> ), .B(n103), .C(n84), .D(n49), .Y(n680) );
  AOI22X1 U709 ( .A(\In<10> ), .B(n16), .C(\In<11> ), .D(n3), .Y(n679) );
  OAI21X1 U710 ( .A(n682), .B(n681), .C(n399), .Y(n688) );
  AOI21X1 U711 ( .A(\In<1> ), .B(n102), .C(n532), .Y(n684) );
  AOI21X1 U712 ( .A(\In<7> ), .B(n72), .C(n142), .Y(n685) );
  OAI21X1 U713 ( .A(n353), .B(n40), .C(n232), .Y(n687) );
  NAND3X1 U714 ( .A(n603), .B(n736), .C(n735), .Y(n698) );
  AOI21X1 U715 ( .A(\In<5> ), .B(n31), .C(n519), .Y(n690) );
  AOI21X1 U716 ( .A(\In<3> ), .B(n68), .C(n289), .Y(n689) );
  AOI22X1 U717 ( .A(\In<5> ), .B(n42), .C(\In<4> ), .D(n49), .Y(n692) );
  AOI22X1 U718 ( .A(\In<6> ), .B(n621), .C(\In<7> ), .D(n20), .Y(n691) );
  OAI21X1 U719 ( .A(n759), .B(n135), .C(n234), .Y(n697) );
  AND2X2 U720 ( .A(n387), .B(n74), .Y(n693) );
  NAND3X1 U721 ( .A(n550), .B(n579), .C(n693), .Y(n731) );
  AOI22X1 U722 ( .A(\In<1> ), .B(n101), .C(\In<0> ), .D(n610), .Y(n695) );
  AOI22X1 U723 ( .A(\In<2> ), .B(n16), .C(\In<3> ), .D(n72), .Y(n694) );
  OAI21X1 U724 ( .A(n758), .B(n160), .C(n236), .Y(n696) );
  NAND3X1 U725 ( .A(n271), .B(n275), .C(n266), .Y(\Out<3> ) );
  OAI21X1 U726 ( .A(n153), .B(n135), .C(n404), .Y(n699) );
  AOI21X1 U727 ( .A(n577), .B(n739), .C(n699), .Y(n704) );
  OAI21X1 U728 ( .A(n700), .B(n158), .C(n406), .Y(n703) );
  OAI21X1 U729 ( .A(n353), .B(n108), .C(n39), .Y(n702) );
  OAI21X1 U730 ( .A(n590), .B(n170), .C(n326), .Y(n706) );
  OAI21X1 U731 ( .A(n595), .B(n322), .C(n408), .Y(n705) );
  OAI21X1 U732 ( .A(n65), .B(n121), .C(n410), .Y(n707) );
  AOI21X1 U733 ( .A(n764), .B(n75), .C(n707), .Y(n708) );
  OAI21X1 U734 ( .A(n547), .B(n121), .C(n412), .Y(n710) );
  OAI21X1 U735 ( .A(n590), .B(n35), .C(n414), .Y(n709) );
  OAI21X1 U736 ( .A(n582), .B(n322), .C(n416), .Y(n711) );
  OAI21X1 U737 ( .A(n40), .B(n559), .C(n418), .Y(n767) );
  AOI21X1 U738 ( .A(n763), .B(n767), .C(n467), .Y(n714) );
  AOI22X1 U739 ( .A(n190), .B(n757), .C(n267), .D(n578), .Y(n713) );
  OAI21X1 U740 ( .A(n43), .B(n149), .C(n360), .Y(n712) );
  NAND3X1 U741 ( .A(n476), .B(n491), .C(n503), .Y(n773) );
  AOI22X1 U742 ( .A(n154), .B(n757), .C(n98), .D(n267), .Y(n719) );
  OAI21X1 U743 ( .A(n322), .B(n716), .C(n419), .Y(n718) );
  OAI21X1 U744 ( .A(n121), .B(n158), .C(n422), .Y(n717) );
  OAI21X1 U745 ( .A(n590), .B(n22), .C(n335), .Y(n720) );
  AOI21X1 U746 ( .A(n575), .B(n764), .C(n720), .Y(n724) );
  AND2X2 U747 ( .A(n144), .B(n48), .Y(n721) );
  AOI21X1 U748 ( .A(n37), .B(n757), .C(n721), .Y(n723) );
  OAI21X1 U749 ( .A(n749), .B(n135), .C(n423), .Y(n722) );
  NAND3X1 U750 ( .A(n493), .B(n52), .C(n477), .Y(\Out<9> ) );
  AOI22X1 U751 ( .A(n726), .B(n548), .C(n739), .D(n573), .Y(n730) );
  AOI22X1 U752 ( .A(n763), .B(n33), .C(n764), .D(n571), .Y(n729) );
  OAI21X1 U753 ( .A(n590), .B(n17), .C(n336), .Y(n728) );
  OAI21X1 U754 ( .A(n353), .B(n528), .C(n424), .Y(n727) );
  NAND3X1 U755 ( .A(n471), .B(n492), .C(n505), .Y(\Out<10> ) );
  AND2X2 U756 ( .A(n768), .B(n557), .Y(n732) );
  AOI22X1 U757 ( .A(n570), .B(n732), .C(n739), .D(n552), .Y(n738) );
  NAND3X1 U758 ( .A(n479), .B(n495), .C(n506), .Y(n734) );
  NAND3X1 U759 ( .A(n344), .B(n346), .C(n508), .Y(n733) );
  NAND3X1 U760 ( .A(n736), .B(n735), .C(n600), .Y(n737) );
  AOI22X1 U761 ( .A(n117), .B(n739), .C(n27), .D(n267), .Y(n746) );
  AND2X2 U762 ( .A(n740), .B(n603), .Y(n743) );
  OAI21X1 U763 ( .A(n158), .B(n135), .C(n368), .Y(n742) );
  OAI21X1 U764 ( .A(n143), .B(n153), .C(n425), .Y(n745) );
  NAND3X1 U765 ( .A(n472), .B(n58), .C(n56), .Y(\Out<12> ) );
  OAI21X1 U766 ( .A(n562), .B(n170), .C(n427), .Y(n748) );
  OAI21X1 U767 ( .A(n83), .B(n595), .C(n371), .Y(n747) );
  OAI21X1 U768 ( .A(n353), .B(n65), .C(n374), .Y(n750) );
  AOI21X1 U769 ( .A(n762), .B(n75), .C(n750), .Y(n752) );
  NAND3X1 U770 ( .A(n15), .B(n498), .C(n500), .Y(n772) );
  OAI21X1 U771 ( .A(n83), .B(n582), .C(n429), .Y(n755) );
  OAI21X1 U772 ( .A(n562), .B(n35), .C(n376), .Y(n754) );
  OAI21X1 U773 ( .A(n353), .B(n547), .C(n430), .Y(n756) );
  OAI21X1 U774 ( .A(n590), .B(n43), .C(n329), .Y(n761) );
  OAI21X1 U775 ( .A(n546), .B(n759), .C(n380), .Y(n760) );
  AOI22X1 U776 ( .A(n763), .B(n578), .C(n762), .D(n93), .Y(n765) );
  AOI21X1 U777 ( .A(n483), .B(n481), .C(\Op<1> ), .Y(n766) );
endmodule


module CLA16_0 ( .A({\A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , 
        \A<9> , \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , 
        \A<0> }), .B({\B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , 
        \B<9> , \B<8> , \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , 
        \B<0> }), Cin, Cout, .S({\S<15> , \S<14> , \S<13> , \S<12> , \S<11> , 
        \S<10> , \S<9> , \S<8> , \S<7> , \S<6> , \S<5> , \S<4> , \S<3> , 
        \S<2> , \S<1> , \S<0> }) );
  input \A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> , \A<8> ,
         \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , \A<0> ,
         \B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , \B<9> , \B<8> ,
         \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output Cout, \S<15> , \S<14> , \S<13> , \S<12> , \S<11> , \S<10> , \S<9> ,
         \S<8> , \S<7> , \S<6> , \S<5> , \S<4> , \S<3> , \S<2> , \S<1> ,
         \S<0> ;
  wire   p30, g30, p74, g74, p118, g118, p1512, g1512, n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33;

  CLA4_3 A3_0 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), .Cin(Cin), .Cout(), .P(p30), .G(g30), .S({\S<3> , 
        \S<2> , \S<1> , \S<0> }) );
  CLA4_2 A7_4 ( .A({\A<7> , \A<6> , \A<5> , \A<4> }), .B({\B<7> , \B<6> , 
        \B<5> , \B<4> }), .Cin(n33), .Cout(), .P(p74), .G(g74), .S({\S<7> , 
        \S<6> , \S<5> , \S<4> }) );
  CLA4_1 A11_8 ( .A({\A<11> , \A<10> , \A<9> , \A<8> }), .B({\B<11> , \B<10> , 
        \B<9> , n9}), .Cin(n30), .Cout(), .P(p118), .G(g118), .S({\S<11> , 
        \S<10> , \S<9> , \S<8> }) );
  CLA4_0 A15_12 ( .A({\A<15> , \A<14> , \A<13> , \A<12> }), .B({\B<15> , 
        \B<14> , \B<13> , \B<12> }), .Cin(n31), .Cout(), .P(p1512), .G(g1512), 
        .S({\S<15> , \S<14> , \S<13> , \S<12> }) );
  INVX1 U1 ( .A(g30), .Y(n1) );
  INVX1 U2 ( .A(g1512), .Y(n27) );
  BUFX2 U3 ( .A(p30), .Y(n2) );
  INVX4 U4 ( .A(n17), .Y(n30) );
  INVX1 U5 ( .A(g30), .Y(n3) );
  INVX1 U6 ( .A(n30), .Y(n4) );
  INVX1 U7 ( .A(n4), .Y(n5) );
  BUFX2 U8 ( .A(p74), .Y(n6) );
  INVX1 U9 ( .A(p118), .Y(n7) );
  INVX1 U10 ( .A(\B<8> ), .Y(n8) );
  INVX1 U11 ( .A(n8), .Y(n9) );
  INVX1 U12 ( .A(g74), .Y(n25) );
  INVX4 U13 ( .A(n20), .Y(n33) );
  AND2X2 U14 ( .A(p30), .B(Cin), .Y(n10) );
  INVX1 U15 ( .A(n10), .Y(n11) );
  BUFX2 U16 ( .A(n26), .Y(n12) );
  BUFX2 U17 ( .A(n29), .Y(n13) );
  OR2X2 U18 ( .A(g74), .B(g118), .Y(n14) );
  INVX1 U19 ( .A(n14), .Y(n15) );
  INVX1 U20 ( .A(n10), .Y(n16) );
  AND2X2 U21 ( .A(n12), .B(n25), .Y(n17) );
  INVX1 U22 ( .A(p1512), .Y(n28) );
  INVX1 U23 ( .A(n3), .Y(n18) );
  INVX1 U24 ( .A(g118), .Y(n23) );
  INVX1 U25 ( .A(n11), .Y(n24) );
  INVX1 U26 ( .A(n23), .Y(n19) );
  AND2X2 U27 ( .A(n16), .B(n1), .Y(n20) );
  AND2X2 U28 ( .A(n2), .B(Cin), .Y(n21) );
  OAI21X1 U29 ( .A(n18), .B(n21), .C(n6), .Y(n22) );
  AOI22X1 U30 ( .A(n23), .B(n7), .C(n22), .D(n15), .Y(n31) );
  AOI22X1 U31 ( .A(g30), .B(p74), .C(p74), .D(n24), .Y(n26) );
  AOI21X1 U32 ( .A(n5), .B(p118), .C(n19), .Y(n29) );
  OAI21X1 U33 ( .A(n13), .B(n28), .C(n27), .Y(Cout) );
endmodule


module dff_451 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_450 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_449 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_448 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_447 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_446 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_445 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_444 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_443 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_442 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_441 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_440 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_439 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_438 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_437 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_436 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_435 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_434 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_433 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_432 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_431 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_430 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_429 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_428 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_427 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_426 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_425 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_424 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_423 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_422 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_421 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_420 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_419 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_418 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_417 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_416 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_415 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_414 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_413 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_412 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_411 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_410 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_409 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_408 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_407 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_406 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_405 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_404 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_403 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_402 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_401 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_400 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_399 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_398 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_397 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_396 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_395 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_394 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_393 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_392 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_391 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_390 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_389 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_388 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_387 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_386 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_385 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_384 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_383 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_382 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_381 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_380 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_379 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_378 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_377 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_376 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_375 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_374 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_373 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_372 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_371 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_370 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_369 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_368 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_367 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_366 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_365 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_364 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_363 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_362 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_361 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_360 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_359 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_358 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_357 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_356 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_355 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_354 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_353 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_352 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_351 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_350 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_349 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_348 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_347 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_346 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_345 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_344 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_343 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_342 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_341 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_340 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_339 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_338 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_337 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_336 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_335 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_334 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_333 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_332 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_331 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_330 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_329 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX2 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_328 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_327 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_326 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X2 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module dff_325 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_324 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_323 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_322 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_321 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_320 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_319 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_318 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_317 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_316 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_315 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_314 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_313 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_312 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_311 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_310 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_309 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_308 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_307 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_306 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_305 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_304 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_303 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_302 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_301 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_300 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_299 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_298 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_297 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_296 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_295 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_294 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_293 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_292 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_291 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_290 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_289 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_288 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_287 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_286 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_285 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_284 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_283 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_282 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_281 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_280 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_279 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_278 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_277 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_276 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_275 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_274 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_273 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_272 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_271 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_270 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_269 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_268 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_267 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_266 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_265 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_264 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_263 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_262 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_261 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_260 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_259 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_258 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_257 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_256 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_255 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_254 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_253 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_252 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_251 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_250 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_249 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_248 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_247 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_246 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_245 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_244 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_243 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_242 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_241 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_240 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_239 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_238 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_237 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_236 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_235 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_234 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_233 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_232 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_231 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_230 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_229 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_228 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_227 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_226 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_225 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_224 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_223 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_222 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_221 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_220 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_219 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_218 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_217 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_216 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_215 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_214 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_213 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_212 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_211 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_210 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_209 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_208 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_207 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_206 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_205 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_204 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_203 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_202 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_201 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_200 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_199 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_198 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_197 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_196 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_195 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_194 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_193 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_192 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_191 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_190 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_189 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_188 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_187 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_186 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_185 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_184 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_183 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_182 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_181 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_180 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_179 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X1 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_178 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_177 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_176 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_175 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_174 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_173 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_172 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_171 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_170 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_169 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_168 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_167 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_166 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_165 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_164 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_163 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(rst), .B(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n4) );
endmodule


module dff_162 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X2 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_161 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X2 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_160 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n3, n4;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n4) );
  OR2X2 U4 ( .A(rst), .B(n4), .Y(n1) );
  INVX2 U5 ( .A(n1), .Y(n3) );
endmodule


module dff_665 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n2, n1, n3;

  DFFPOSX1 state_reg ( .D(n3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n2) );
  OR2X1 U4 ( .A(rst), .B(n2), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n3) );
endmodule


module reg1_26 ( d, q, clk, rst, en );
  input d, clk, rst, en;
  output q;
  wire   n2, n3, n4, n1;

  dff_664 d0 ( .q(q), .d(n2), .clk(clk), .rst(rst) );
  AOI22X1 U3 ( .A(en), .B(d), .C(q), .D(n3), .Y(n4) );
  INVX1 U1 ( .A(en), .Y(n3) );
  BUFX2 U2 ( .A(n4), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n2) );
endmodule


module reg16_36 ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n1, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49;

  dff_663 d0 ( .q(\read<0> ), .d(n2), .clk(clk), .rst(rst) );
  dff_662 d1 ( .q(\read<1> ), .d(n3), .clk(clk), .rst(rst) );
  dff_661 d2 ( .q(\read<2> ), .d(n4), .clk(clk), .rst(rst) );
  dff_660 d3 ( .q(\read<3> ), .d(n5), .clk(clk), .rst(rst) );
  dff_659 d4 ( .q(\read<4> ), .d(n6), .clk(clk), .rst(rst) );
  dff_658 d5 ( .q(\read<5> ), .d(n7), .clk(clk), .rst(rst) );
  dff_657 d6 ( .q(\read<6> ), .d(n8), .clk(clk), .rst(rst) );
  dff_656 d7 ( .q(\read<7> ), .d(n9), .clk(clk), .rst(rst) );
  dff_655 d8 ( .q(\read<8> ), .d(n10), .clk(clk), .rst(rst) );
  dff_654 d9 ( .q(\read<9> ), .d(n11), .clk(clk), .rst(rst) );
  dff_653 d10 ( .q(\read<10> ), .d(n12), .clk(clk), .rst(rst) );
  dff_652 d11 ( .q(\read<11> ), .d(n13), .clk(clk), .rst(rst) );
  dff_651 d12 ( .q(\read<12> ), .d(n14), .clk(clk), .rst(rst) );
  dff_650 d13 ( .q(\read<13> ), .d(n15), .clk(clk), .rst(rst) );
  dff_649 d14 ( .q(\read<14> ), .d(n16), .clk(clk), .rst(rst) );
  dff_648 d15 ( .q(\read<15> ), .d(n17), .clk(clk), .rst(rst) );
  AOI22X1 U18 ( .A(\read<9> ), .B(n18), .C(\write<9> ), .D(wr_en), .Y(n19) );
  AOI22X1 U19 ( .A(\read<8> ), .B(n18), .C(\write<8> ), .D(wr_en), .Y(n20) );
  AOI22X1 U20 ( .A(\read<7> ), .B(n18), .C(\write<7> ), .D(wr_en), .Y(n21) );
  AOI22X1 U21 ( .A(\read<6> ), .B(n18), .C(\write<6> ), .D(wr_en), .Y(n22) );
  AOI22X1 U22 ( .A(\read<5> ), .B(n18), .C(\write<5> ), .D(wr_en), .Y(n23) );
  AOI22X1 U23 ( .A(\read<4> ), .B(n18), .C(\write<4> ), .D(wr_en), .Y(n24) );
  AOI22X1 U24 ( .A(\read<3> ), .B(n18), .C(\write<3> ), .D(wr_en), .Y(n25) );
  AOI22X1 U25 ( .A(\read<2> ), .B(n18), .C(\write<2> ), .D(wr_en), .Y(n26) );
  AOI22X1 U26 ( .A(\read<1> ), .B(n18), .C(\write<1> ), .D(wr_en), .Y(n27) );
  AOI22X1 U27 ( .A(\read<15> ), .B(n18), .C(\write<15> ), .D(wr_en), .Y(n28)
         );
  AOI22X1 U28 ( .A(\read<14> ), .B(n18), .C(\write<14> ), .D(wr_en), .Y(n29)
         );
  AOI22X1 U29 ( .A(\read<13> ), .B(n18), .C(\write<13> ), .D(wr_en), .Y(n30)
         );
  AOI22X1 U30 ( .A(\read<12> ), .B(n18), .C(\write<12> ), .D(wr_en), .Y(n31)
         );
  AOI22X1 U31 ( .A(\read<11> ), .B(n18), .C(\write<11> ), .D(wr_en), .Y(n32)
         );
  AOI22X1 U32 ( .A(\read<10> ), .B(n18), .C(\write<10> ), .D(wr_en), .Y(n33)
         );
  AOI22X1 U33 ( .A(\read<0> ), .B(n18), .C(\write<0> ), .D(wr_en), .Y(n34) );
  INVX1 U1 ( .A(n1), .Y(n2) );
  INVX1 U2 ( .A(n41), .Y(n3) );
  INVX1 U3 ( .A(n42), .Y(n4) );
  INVX1 U4 ( .A(n43), .Y(n5) );
  INVX1 U5 ( .A(n44), .Y(n6) );
  INVX1 U6 ( .A(n45), .Y(n7) );
  INVX1 U7 ( .A(n46), .Y(n8) );
  INVX1 U8 ( .A(n47), .Y(n9) );
  INVX1 U9 ( .A(n48), .Y(n10) );
  INVX1 U10 ( .A(n49), .Y(n11) );
  INVX1 U11 ( .A(n35), .Y(n12) );
  INVX1 U12 ( .A(n37), .Y(n14) );
  INVX1 U13 ( .A(n38), .Y(n15) );
  INVX1 U14 ( .A(n39), .Y(n16) );
  INVX1 U15 ( .A(n40), .Y(n17) );
  INVX1 U16 ( .A(wr_en), .Y(n18) );
  BUFX2 U17 ( .A(n34), .Y(n1) );
  BUFX2 U34 ( .A(n33), .Y(n35) );
  BUFX2 U35 ( .A(n32), .Y(n36) );
  INVX1 U36 ( .A(n36), .Y(n13) );
  BUFX2 U37 ( .A(n31), .Y(n37) );
  BUFX2 U38 ( .A(n30), .Y(n38) );
  BUFX2 U39 ( .A(n29), .Y(n39) );
  BUFX2 U40 ( .A(n28), .Y(n40) );
  BUFX2 U41 ( .A(n27), .Y(n41) );
  BUFX2 U42 ( .A(n26), .Y(n42) );
  BUFX2 U43 ( .A(n25), .Y(n43) );
  BUFX2 U44 ( .A(n24), .Y(n44) );
  BUFX2 U45 ( .A(n23), .Y(n45) );
  BUFX2 U46 ( .A(n22), .Y(n46) );
  BUFX2 U47 ( .A(n21), .Y(n47) );
  BUFX2 U48 ( .A(n20), .Y(n48) );
  BUFX2 U49 ( .A(n19), .Y(n49) );
endmodule


module IF_control ( Jump, Branch, jmp_r, .opcode({\opcode<4> , \opcode<3> , 
        \opcode<2> , \opcode<1> , \opcode<0> }) );
  input \opcode<4> , \opcode<3> , \opcode<2> , \opcode<1> , \opcode<0> ;
  output Jump, Branch, jmp_r;
  wire   n1, n2;

  NOR3X1 U4 ( .A(\opcode<3> ), .B(\opcode<4> ), .C(n2), .Y(Jump) );
  NOR3X1 U5 ( .A(n1), .B(\opcode<4> ), .C(n2), .Y(Branch) );
  INVX1 U1 ( .A(\opcode<3> ), .Y(n1) );
  INVX1 U2 ( .A(\opcode<2> ), .Y(n2) );
  AND2X1 U3 ( .A(\opcode<0> ), .B(Jump), .Y(jmp_r) );
endmodule


module pc ( branch_if, .pc_inc_two({\pc_inc_two<15> , \pc_inc_two<14> , 
        \pc_inc_two<13> , \pc_inc_two<12> , \pc_inc_two<11> , \pc_inc_two<10> , 
        \pc_inc_two<9> , \pc_inc_two<8> , \pc_inc_two<7> , \pc_inc_two<6> , 
        \pc_inc_two<5> , \pc_inc_two<4> , \pc_inc_two<3> , \pc_inc_two<2> , 
        \pc_inc_two<1> , \pc_inc_two<0> }), jmp_r, en, clk, rst, jump, .inst({
        \inst<15> , \inst<14> , \inst<13> , \inst<12> , \inst<11> , \inst<10> , 
        \inst<9> , \inst<8> , \inst<7> , \inst<6> , \inst<5> , \inst<4> , 
        \inst<3> , \inst<2> , \inst<1> , \inst<0> }), .addr({\addr<15> , 
        \addr<14> , \addr<13> , \addr<12> , \addr<11> , \addr<10> , \addr<9> , 
        \addr<8> , \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , 
        \addr<2> , \addr<1> , \addr<0> }), branch, .rs({\rs<15> , \rs<14> , 
        \rs<13> , \rs<12> , \rs<11> , \rs<10> , \rs<9> , \rs<8> , \rs<7> , 
        \rs<6> , \rs<5> , \rs<4> , \rs<3> , \rs<2> , \rs<1> , \rs<0> }), 
    .pc_nx({\pc_nx<15> , \pc_nx<14> , \pc_nx<13> , \pc_nx<12> , \pc_nx<11> , 
        \pc_nx<10> , \pc_nx<9> , \pc_nx<8> , \pc_nx<7> , \pc_nx<6> , 
        \pc_nx<5> , \pc_nx<4> , \pc_nx<3> , \pc_nx<2> , \pc_nx<1> , \pc_nx<0> 
        }), .EX_inst({\EX_inst<15> , \EX_inst<14> , \EX_inst<13> , 
        \EX_inst<12> , \EX_inst<11> , \EX_inst<10> , \EX_inst<9> , 
        \EX_inst<8> , \EX_inst<7> , \EX_inst<6> , \EX_inst<5> , \EX_inst<4> , 
        \EX_inst<3> , \EX_inst<2> , \EX_inst<1> , \EX_inst<0> }), br_ctl );
  input branch_if, jmp_r, en, clk, rst, jump, \inst<15> , \inst<14> ,
         \inst<13> , \inst<12> , \inst<11> , \inst<10> , \inst<9> , \inst<8> ,
         \inst<7> , \inst<6> , \inst<5> , \inst<4> , \inst<3> , \inst<2> ,
         \inst<1> , \inst<0> , branch, \rs<15> , \rs<14> , \rs<13> , \rs<12> ,
         \rs<11> , \rs<10> , \rs<9> , \rs<8> , \rs<7> , \rs<6> , \rs<5> ,
         \rs<4> , \rs<3> , \rs<2> , \rs<1> , \rs<0> , \EX_inst<15> ,
         \EX_inst<14> , \EX_inst<13> , \EX_inst<12> , \EX_inst<11> ,
         \EX_inst<10> , \EX_inst<9> , \EX_inst<8> , \EX_inst<7> , \EX_inst<6> ,
         \EX_inst<5> , \EX_inst<4> , \EX_inst<3> , \EX_inst<2> , \EX_inst<1> ,
         \EX_inst<0> ;
  output \pc_inc_two<15> , \pc_inc_two<14> , \pc_inc_two<13> ,
         \pc_inc_two<12> , \pc_inc_two<11> , \pc_inc_two<10> , \pc_inc_two<9> ,
         \pc_inc_two<8> , \pc_inc_two<7> , \pc_inc_two<6> , \pc_inc_two<5> ,
         \pc_inc_two<4> , \pc_inc_two<3> , \pc_inc_two<2> , \pc_inc_two<1> ,
         \pc_inc_two<0> , \addr<15> , \addr<14> , \addr<13> , \addr<12> ,
         \addr<11> , \addr<10> , \addr<9> , \addr<8> , \addr<7> , \addr<6> ,
         \addr<5> , \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> ,
         \pc_nx<15> , \pc_nx<14> , \pc_nx<13> , \pc_nx<12> , \pc_nx<11> ,
         \pc_nx<10> , \pc_nx<9> , \pc_nx<8> , \pc_nx<7> , \pc_nx<6> ,
         \pc_nx<5> , \pc_nx<4> , \pc_nx<3> , \pc_nx<2> , \pc_nx<1> ,
         \pc_nx<0> , br_ctl;
  wire   n199, n200, n201, n202, n203, n204, n205, n206, n207,
         \branch_addr<15> , \branch_addr<14> , \branch_addr<13> ,
         \branch_addr<12> , \branch_addr<11> , \branch_addr<10> ,
         \branch_addr<9> , \branch_addr<8> , \branch_addr<7> ,
         \branch_addr<6> , \branch_addr<5> , \branch_addr<4> ,
         \branch_addr<3> , \branch_addr<2> , \branch_addr<1> ,
         \branch_addr<0> , \br_inc<15> , \br_inc<14> , \br_inc<13> ,
         \br_inc<12> , \br_inc<11> , \br_inc<10> , \br_inc<9> , \br_inc<8> ,
         \br_inc<7> , \br_inc<6> , \br_inc<5> , \br_inc<4> , \br_inc<3> ,
         \br_inc<2> , \br_inc<1> , \br_inc<0> , \br_pre<15> , \br_pre<14> ,
         \br_pre<13> , \br_pre<12> , \br_pre<11> , \br_pre<10> , \br_pre<9> ,
         \br_pre<8> , \br_pre<7> , \br_pre<6> , \br_pre<5> , \br_pre<4> ,
         \br_pre<3> , \br_pre<2> , \br_pre<1> , \br_pre<0> , \jmp_d<15> ,
         \jmp_d<14> , \jmp_d<13> , \jmp_d<12> , \jmp_d<11> , \jmp_d<10> ,
         \jmp_d<9> , \jmp_d<8> , \jmp_d<7> , \jmp_d<6> , \jmp_d<5> ,
         \jmp_d<4> , \jmp_d<3> , \jmp_d<2> , \jmp_d<1> , \jmp_d<0> ,
         \jmp_i<15> , \jmp_i<14> , \jmp_i<13> , \jmp_i<12> , \jmp_i<11> ,
         \jmp_i<10> , \jmp_i<9> , \jmp_i<8> , \jmp_i<7> , \jmp_i<6> ,
         \jmp_i<5> , \jmp_i<4> , \jmp_i<3> , \jmp_i<2> , \jmp_i<1> ,
         \jmp_i<0> , n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n60, n63, n65, n66, n68, n69, n70, n72, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n126, n128, n130,
         n132, n135, n136, n137, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198;

  reg16_9 branch_addr_reg ( .read({\branch_addr<15> , \branch_addr<14> , 
        \branch_addr<13> , \branch_addr<12> , \branch_addr<11> , 
        \branch_addr<10> , \branch_addr<9> , \branch_addr<8> , 
        \branch_addr<7> , \branch_addr<6> , \branch_addr<5> , \branch_addr<4> , 
        \branch_addr<3> , \branch_addr<2> , \branch_addr<1> , \branch_addr<0> }), .write({\addr<15> , \addr<14> , \addr<13> , \addr<12> , \addr<11> , 
        \addr<10> , \addr<9> , \addr<8> , \addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , n3, \addr<1> , \addr<0> }), .wr_en(branch_if), 
        .rst(rst), .clk(clk) );
  reg16_8 pc_dff ( .read({\addr<15> , \addr<14> , \addr<13> , \addr<12> , 
        \addr<11> , \addr<10> , \addr<9> , \addr<8> , \addr<7> , \addr<6> , 
        \addr<5> , \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), 
        .write({n198, \pc_nx<14> , \pc_nx<13> , n141, \pc_nx<11> , n136, 
        \pc_nx<9> , n70, \pc_nx<7> , \pc_nx<6> , n68, \pc_nx<4> , \pc_nx<3> , 
        \pc_nx<2> , \pc_nx<1> , n65}), .wr_en(en), .rst(rst), .clk(clk) );
  CLA16_5 pc_incr ( .A({\addr<15> , \addr<14> , \addr<13> , \addr<12> , 
        \addr<11> , \addr<10> , \addr<9> , \addr<8> , \addr<7> , \addr<6> , 
        \addr<5> , \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b1, 1'b0}), .Cin(1'b0), .Cout(), .S({
        \pc_inc_two<15> , \pc_inc_two<14> , \pc_inc_two<13> , \pc_inc_two<12> , 
        n199, \pc_inc_two<10> , \pc_inc_two<9> , \pc_inc_two<8> , n200, n201, 
        n202, \pc_inc_two<4> , \pc_inc_two<3> , \pc_inc_two<2> , 
        \pc_inc_two<1> , \pc_inc_two<0> }) );
  CLA16_4 br_inc_two ( .A({\branch_addr<15> , \branch_addr<14> , 
        \branch_addr<13> , \branch_addr<12> , \branch_addr<11> , 
        \branch_addr<10> , \branch_addr<9> , \branch_addr<8> , 
        \branch_addr<7> , \branch_addr<6> , \branch_addr<5> , \branch_addr<4> , 
        \branch_addr<3> , \branch_addr<2> , \branch_addr<1> , \branch_addr<0> }), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b1, 1'b0}), .Cin(1'b0), .Cout(), .S({\br_inc<15> , 
        \br_inc<14> , \br_inc<13> , \br_inc<12> , \br_inc<11> , \br_inc<10> , 
        \br_inc<9> , \br_inc<8> , \br_inc<7> , \br_inc<6> , \br_inc<5> , 
        \br_inc<4> , \br_inc<3> , \br_inc<2> , \br_inc<1> , \br_inc<0> }) );
  CLA16_3 br_add ( .A({\br_inc<15> , \br_inc<14> , \br_inc<13> , \br_inc<12> , 
        \br_inc<11> , \br_inc<10> , \br_inc<9> , \br_inc<8> , \br_inc<7> , 
        \br_inc<6> , \br_inc<5> , \br_inc<4> , \br_inc<3> , \br_inc<2> , 
        \br_inc<1> , \br_inc<0> }), .B({n163, n163, n163, n164, n164, n164, 
        n164, n164, n164, \EX_inst<6> , \EX_inst<5> , \EX_inst<4> , 
        \EX_inst<3> , \EX_inst<2> , \EX_inst<1> , \EX_inst<0> }), .Cin(1'b0), 
        .Cout(), .S({\br_pre<15> , \br_pre<14> , \br_pre<13> , \br_pre<12> , 
        \br_pre<11> , \br_pre<10> , \br_pre<9> , \br_pre<8> , \br_pre<7> , 
        \br_pre<6> , \br_pre<5> , \br_pre<4> , \br_pre<3> , \br_pre<2> , 
        \br_pre<1> , \br_pre<0> }) );
  CLA16_2 jmp_add_d ( .A({\pc_inc_two<15> , \pc_inc_two<14> , \pc_inc_two<13> , 
        \pc_inc_two<12> , n199, \pc_inc_two<10> , \pc_inc_two<9> , 
        \pc_inc_two<8> , n200, n201, n202, \pc_inc_two<4> , \pc_inc_two<3> , 
        \pc_inc_two<2> , \pc_inc_two<1> , \pc_inc_two<0> }), .B({\EX_inst<10> , 
        \EX_inst<10> , \EX_inst<10> , \EX_inst<10> , \EX_inst<10> , 
        \EX_inst<10> , \EX_inst<9> , \EX_inst<8> , n163, \EX_inst<6> , 
        \EX_inst<5> , \EX_inst<4> , \EX_inst<3> , \EX_inst<2> , \EX_inst<1> , 
        \EX_inst<0> }), .Cin(1'b0), .Cout(), .S({\jmp_d<15> , \jmp_d<14> , 
        \jmp_d<13> , \jmp_d<12> , \jmp_d<11> , \jmp_d<10> , \jmp_d<9> , 
        \jmp_d<8> , \jmp_d<7> , \jmp_d<6> , \jmp_d<5> , \jmp_d<4> , \jmp_d<3> , 
        \jmp_d<2> , \jmp_d<1> , \jmp_d<0> }) );
  CLA16_1 jmp_add_i ( .A({\rs<15> , n148, n77, \rs<12> , n157, n85, n79, n153, 
        \rs<7> , n80, \rs<5> , n78, n86, n150, \rs<1> , \rs<0> }), .B({n163, 
        n163, n163, n163, n163, n163, n163, n163, n163, \EX_inst<6> , 
        \EX_inst<5> , \EX_inst<4> , \EX_inst<3> , \EX_inst<2> , \EX_inst<1> , 
        \EX_inst<0> }), .Cin(1'b0), .Cout(), .S({\jmp_i<15> , \jmp_i<14> , 
        \jmp_i<13> , \jmp_i<12> , \jmp_i<11> , \jmp_i<10> , \jmp_i<9> , 
        \jmp_i<8> , \jmp_i<7> , \jmp_i<6> , \jmp_i<5> , \jmp_i<4> , \jmp_i<3> , 
        \jmp_i<2> , \jmp_i<1> , \jmp_i<0> }) );
  AND2X2 U3 ( .A(n93), .B(n100), .Y(n135) );
  AND2X2 U4 ( .A(n16), .B(n25), .Y(n72) );
  INVX1 U5 ( .A(n165), .Y(n164) );
  INVX1 U6 ( .A(\EX_inst<7> ), .Y(n165) );
  AND2X1 U7 ( .A(n20), .B(n31), .Y(n40) );
  AND2X1 U8 ( .A(\EX_inst<14> ), .B(\EX_inst<13> ), .Y(n160) );
  OR2X1 U9 ( .A(n169), .B(\EX_inst<15> ), .Y(n34) );
  INVX1 U10 ( .A(jump), .Y(n171) );
  AND2X1 U11 ( .A(jump), .B(\EX_inst<11> ), .Y(n122) );
  AND2X1 U12 ( .A(n10), .B(n37), .Y(n4) );
  AND2X1 U13 ( .A(\jmp_i<11> ), .B(n122), .Y(n90) );
  BUFX2 U14 ( .A(n202), .Y(\pc_inc_two<5> ) );
  AND2X2 U15 ( .A(\br_pre<15> ), .B(n195), .Y(n144) );
  BUFX2 U16 ( .A(\rs<4> ), .Y(n78) );
  AND2X2 U17 ( .A(\br_pre<14> ), .B(n195), .Y(n105) );
  BUFX2 U18 ( .A(n201), .Y(\pc_inc_two<6> ) );
  BUFX2 U19 ( .A(\addr<2> ), .Y(n3) );
  AND2X1 U20 ( .A(\jmp_i<14> ), .B(n122), .Y(n110) );
  OR2X2 U21 ( .A(n123), .B(n91), .Y(n88) );
  OR2X2 U22 ( .A(n90), .B(n88), .Y(\pc_nx<11> ) );
  INVX1 U23 ( .A(\EX_inst<11> ), .Y(n161) );
  OR2X2 U24 ( .A(n79), .B(\rs<8> ), .Y(n5) );
  INVX1 U25 ( .A(n5), .Y(n6) );
  AND2X2 U26 ( .A(\rs<15> ), .B(\EX_inst<11> ), .Y(n7) );
  INVX1 U27 ( .A(n7), .Y(n8) );
  AND2X2 U28 ( .A(\br_pre<0> ), .B(n195), .Y(n9) );
  INVX1 U29 ( .A(n9), .Y(n10) );
  AND2X2 U30 ( .A(n171), .B(n60), .Y(n11) );
  INVX1 U31 ( .A(n11), .Y(n12) );
  AND2X2 U32 ( .A(\pc_inc_two<2> ), .B(n196), .Y(n13) );
  INVX1 U33 ( .A(n13), .Y(n14) );
  BUFX2 U34 ( .A(n184), .Y(n15) );
  BUFX2 U35 ( .A(n186), .Y(n16) );
  OR2X2 U36 ( .A(\rs<15> ), .B(\rs<14> ), .Y(n17) );
  INVX1 U37 ( .A(n17), .Y(n18) );
  OR2X2 U38 ( .A(\rs<0> ), .B(n152), .Y(n19) );
  INVX1 U39 ( .A(n19), .Y(n20) );
  OR2X2 U40 ( .A(\rs<7> ), .B(n80), .Y(n21) );
  INVX1 U41 ( .A(n21), .Y(n22) );
  BUFX2 U42 ( .A(n177), .Y(n23) );
  BUFX2 U43 ( .A(n183), .Y(n24) );
  BUFX2 U44 ( .A(n185), .Y(n25) );
  OR2X2 U45 ( .A(n85), .B(\rs<11> ), .Y(n26) );
  INVX1 U46 ( .A(n26), .Y(n27) );
  OR2X2 U47 ( .A(n77), .B(\rs<12> ), .Y(n28) );
  INVX1 U48 ( .A(n28), .Y(n29) );
  OR2X2 U49 ( .A(n150), .B(n86), .Y(n30) );
  INVX1 U50 ( .A(n30), .Y(n31) );
  OR2X2 U51 ( .A(n78), .B(\rs<5> ), .Y(n32) );
  INVX1 U52 ( .A(n32), .Y(n33) );
  INVX1 U53 ( .A(n34), .Y(n35) );
  AND2X2 U54 ( .A(\pc_inc_two<0> ), .B(n196), .Y(n36) );
  INVX1 U55 ( .A(n36), .Y(n37) );
  AND2X2 U56 ( .A(n18), .B(n29), .Y(n38) );
  INVX1 U57 ( .A(n38), .Y(n39) );
  INVX1 U58 ( .A(n40), .Y(n41) );
  AND2X2 U59 ( .A(n6), .B(n27), .Y(n42) );
  INVX1 U60 ( .A(n42), .Y(n43) );
  AND2X2 U61 ( .A(n22), .B(n33), .Y(n44) );
  INVX1 U62 ( .A(n44), .Y(n45) );
  AND2X2 U63 ( .A(\br_pre<1> ), .B(n195), .Y(n46) );
  INVX1 U64 ( .A(n46), .Y(n47) );
  AND2X2 U65 ( .A(\br_pre<2> ), .B(n195), .Y(n48) );
  INVX1 U66 ( .A(n48), .Y(n49) );
  AND2X2 U67 ( .A(\br_pre<3> ), .B(n195), .Y(n50) );
  INVX1 U68 ( .A(n50), .Y(n51) );
  AND2X2 U69 ( .A(\br_pre<4> ), .B(n195), .Y(n52) );
  INVX1 U70 ( .A(n52), .Y(n53) );
  AND2X2 U71 ( .A(n82), .B(n147), .Y(n54) );
  INVX1 U72 ( .A(n54), .Y(n55) );
  BUFX2 U73 ( .A(n175), .Y(n56) );
  AND2X2 U74 ( .A(\pc_inc_two<1> ), .B(n196), .Y(n57) );
  INVX1 U75 ( .A(n57), .Y(n58) );
  AND2X2 U76 ( .A(n170), .B(n35), .Y(br_ctl) );
  INVX1 U77 ( .A(br_ctl), .Y(n60) );
  BUFX2 U78 ( .A(n204), .Y(\pc_nx<4> ) );
  BUFX2 U79 ( .A(n203), .Y(\pc_nx<14> ) );
  AND2X2 U80 ( .A(n107), .B(n4), .Y(n63) );
  INVX1 U81 ( .A(n63), .Y(\pc_nx<0> ) );
  INVX1 U82 ( .A(n63), .Y(n65) );
  AND2X2 U83 ( .A(n109), .B(n23), .Y(n66) );
  INVX1 U84 ( .A(n66), .Y(\pc_nx<5> ) );
  INVX1 U85 ( .A(n66), .Y(n68) );
  AND2X2 U86 ( .A(n15), .B(n24), .Y(n69) );
  INVX1 U87 ( .A(n69), .Y(n70) );
  INVX1 U88 ( .A(n69), .Y(\pc_nx<8> ) );
  INVX1 U89 ( .A(n72), .Y(\pc_nx<9> ) );
  OR2X2 U90 ( .A(n41), .B(n45), .Y(n74) );
  INVX1 U91 ( .A(n74), .Y(n75) );
  INVX1 U92 ( .A(n74), .Y(n76) );
  BUFX2 U93 ( .A(\rs<13> ), .Y(n77) );
  BUFX2 U94 ( .A(\rs<9> ), .Y(n79) );
  BUFX2 U95 ( .A(\rs<6> ), .Y(n80) );
  OR2X2 U96 ( .A(n39), .B(n43), .Y(n81) );
  INVX1 U97 ( .A(n81), .Y(n82) );
  AND2X2 U98 ( .A(n171), .B(br_ctl), .Y(n83) );
  INVX1 U99 ( .A(n83), .Y(n84) );
  BUFX2 U100 ( .A(\rs<10> ), .Y(n85) );
  BUFX2 U101 ( .A(\rs<3> ), .Y(n86) );
  AND2X1 U102 ( .A(jump), .B(n161), .Y(n89) );
  AND2X1 U103 ( .A(\pc_inc_two<11> ), .B(n196), .Y(n91) );
  BUFX2 U104 ( .A(n180), .Y(n92) );
  BUFX2 U105 ( .A(n182), .Y(n93) );
  BUFX2 U106 ( .A(n188), .Y(n94) );
  BUFX2 U107 ( .A(n191), .Y(n95) );
  BUFX2 U108 ( .A(n193), .Y(n96) );
  AND2X1 U109 ( .A(\jmp_d<14> ), .B(n89), .Y(n97) );
  INVX1 U110 ( .A(n97), .Y(n98) );
  BUFX2 U111 ( .A(n179), .Y(n99) );
  BUFX2 U112 ( .A(n181), .Y(n100) );
  BUFX2 U113 ( .A(n187), .Y(n101) );
  BUFX2 U114 ( .A(n190), .Y(n102) );
  INVX1 U115 ( .A(n192), .Y(n103) );
  INVX1 U116 ( .A(n103), .Y(n104) );
  INVX1 U117 ( .A(n105), .Y(n106) );
  BUFX2 U118 ( .A(n172), .Y(n107) );
  INVX1 U119 ( .A(n178), .Y(n108) );
  INVX1 U120 ( .A(n108), .Y(n109) );
  INVX1 U121 ( .A(n110), .Y(n111) );
  AND2X2 U122 ( .A(\pc_inc_two<3> ), .B(n196), .Y(n112) );
  INVX1 U123 ( .A(n112), .Y(n113) );
  AND2X2 U124 ( .A(\pc_inc_two<4> ), .B(n196), .Y(n114) );
  INVX1 U125 ( .A(n114), .Y(n115) );
  AND2X1 U126 ( .A(\pc_inc_two<14> ), .B(n196), .Y(n116) );
  INVX1 U127 ( .A(n116), .Y(n117) );
  BUFX2 U128 ( .A(n173), .Y(n118) );
  BUFX2 U129 ( .A(n174), .Y(n119) );
  INVX1 U130 ( .A(n176), .Y(n120) );
  INVX1 U131 ( .A(n120), .Y(n121) );
  INVX1 U132 ( .A(n189), .Y(n123) );
  AND2X2 U133 ( .A(n92), .B(n99), .Y(n124) );
  INVX1 U134 ( .A(n124), .Y(\pc_nx<6> ) );
  AND2X2 U135 ( .A(n96), .B(n104), .Y(n126) );
  INVX1 U136 ( .A(n126), .Y(\pc_nx<13> ) );
  INVX1 U137 ( .A(n207), .Y(n128) );
  INVX1 U138 ( .A(n128), .Y(\pc_nx<1> ) );
  INVX1 U139 ( .A(n206), .Y(n130) );
  INVX1 U140 ( .A(n130), .Y(\pc_nx<2> ) );
  INVX1 U141 ( .A(n205), .Y(n132) );
  INVX1 U142 ( .A(n132), .Y(\pc_nx<3> ) );
  INVX1 U143 ( .A(n135), .Y(\pc_nx<7> ) );
  INVX1 U144 ( .A(n137), .Y(n136) );
  AND2X2 U145 ( .A(n94), .B(n101), .Y(n137) );
  INVX1 U146 ( .A(n137), .Y(\pc_nx<10> ) );
  INVX1 U147 ( .A(n140), .Y(\pc_nx<12> ) );
  AND2X2 U148 ( .A(n95), .B(n102), .Y(n140) );
  INVX1 U149 ( .A(n140), .Y(n141) );
  AND2X1 U150 ( .A(\jmp_d<15> ), .B(n89), .Y(n142) );
  INVX1 U151 ( .A(n142), .Y(n143) );
  INVX1 U152 ( .A(n144), .Y(n145) );
  BUFX2 U153 ( .A(n197), .Y(n146) );
  AND2X2 U154 ( .A(n75), .B(n167), .Y(n147) );
  BUFX2 U155 ( .A(\rs<14> ), .Y(n148) );
  INVX1 U156 ( .A(\rs<2> ), .Y(n149) );
  INVX1 U157 ( .A(n149), .Y(n150) );
  INVX1 U158 ( .A(\rs<1> ), .Y(n151) );
  INVX1 U159 ( .A(n151), .Y(n152) );
  BUFX2 U160 ( .A(\rs<8> ), .Y(n153) );
  INVX1 U161 ( .A(\EX_inst<12> ), .Y(n167) );
  BUFX2 U162 ( .A(n200), .Y(\pc_inc_two<7> ) );
  AND2X2 U163 ( .A(n98), .B(n106), .Y(n194) );
  BUFX2 U164 ( .A(n199), .Y(\pc_inc_two<11> ) );
  INVX1 U165 ( .A(\rs<11> ), .Y(n156) );
  INVX1 U166 ( .A(n156), .Y(n157) );
  MUX2X1 U167 ( .B(n168), .A(n55), .S(\EX_inst<11> ), .Y(n169) );
  INVX1 U168 ( .A(n158), .Y(n170) );
  INVX1 U169 ( .A(n166), .Y(n159) );
  OAI21X1 U170 ( .A(n162), .B(n159), .C(n160), .Y(n158) );
  AND2X2 U171 ( .A(n82), .B(n76), .Y(n162) );
  INVX4 U172 ( .A(n84), .Y(n195) );
  INVX4 U173 ( .A(n12), .Y(n196) );
  INVX8 U174 ( .A(n165), .Y(n163) );
  MUX2X1 U175 ( .B(\EX_inst<11> ), .A(n8), .S(\EX_inst<12> ), .Y(n166) );
  OR2X2 U176 ( .A(\rs<15> ), .B(n167), .Y(n168) );
  AOI22X1 U177 ( .A(\jmp_d<0> ), .B(n89), .C(\jmp_i<0> ), .D(n122), .Y(n172)
         );
  AOI22X1 U178 ( .A(\jmp_d<1> ), .B(n89), .C(\jmp_i<1> ), .D(n122), .Y(n173)
         );
  NAND3X1 U179 ( .A(n47), .B(n58), .C(n118), .Y(n207) );
  AOI22X1 U180 ( .A(\jmp_d<2> ), .B(n89), .C(\jmp_i<2> ), .D(n122), .Y(n174)
         );
  NAND3X1 U181 ( .A(n49), .B(n14), .C(n119), .Y(n206) );
  AOI22X1 U182 ( .A(\jmp_d<3> ), .B(n89), .C(\jmp_i<3> ), .D(n122), .Y(n175)
         );
  NAND3X1 U183 ( .A(n51), .B(n56), .C(n113), .Y(n205) );
  AOI22X1 U184 ( .A(\jmp_d<4> ), .B(n89), .C(\jmp_i<4> ), .D(n122), .Y(n176)
         );
  NAND3X1 U185 ( .A(n53), .B(n115), .C(n121), .Y(n204) );
  AOI22X1 U186 ( .A(\jmp_d<5> ), .B(n89), .C(\jmp_i<5> ), .D(n122), .Y(n178)
         );
  AOI22X1 U187 ( .A(\pc_inc_two<5> ), .B(n196), .C(\br_pre<5> ), .D(n195), .Y(
        n177) );
  AOI22X1 U188 ( .A(\jmp_d<6> ), .B(n89), .C(n122), .D(\jmp_i<6> ), .Y(n180)
         );
  AOI22X1 U189 ( .A(\pc_inc_two<6> ), .B(n196), .C(\br_pre<6> ), .D(n195), .Y(
        n179) );
  AOI22X1 U190 ( .A(\jmp_d<7> ), .B(n89), .C(n122), .D(\jmp_i<7> ), .Y(n182)
         );
  AOI22X1 U191 ( .A(\pc_inc_two<7> ), .B(n196), .C(\br_pre<7> ), .D(n195), .Y(
        n181) );
  AOI22X1 U192 ( .A(\jmp_d<8> ), .B(n89), .C(\jmp_i<8> ), .D(n122), .Y(n184)
         );
  AOI22X1 U193 ( .A(\pc_inc_two<8> ), .B(n196), .C(\br_pre<8> ), .D(n195), .Y(
        n183) );
  AOI22X1 U194 ( .A(\jmp_d<9> ), .B(n89), .C(n122), .D(\jmp_i<9> ), .Y(n186)
         );
  AOI22X1 U195 ( .A(\pc_inc_two<9> ), .B(n196), .C(\br_pre<9> ), .D(n195), .Y(
        n185) );
  AOI22X1 U196 ( .A(\jmp_d<10> ), .B(n89), .C(n122), .D(\jmp_i<10> ), .Y(n188)
         );
  AOI22X1 U197 ( .A(\pc_inc_two<10> ), .B(n196), .C(n195), .D(\br_pre<10> ), 
        .Y(n187) );
  AOI22X1 U198 ( .A(n89), .B(\jmp_d<11> ), .C(n195), .D(\br_pre<11> ), .Y(n189) );
  AOI22X1 U199 ( .A(\jmp_d<12> ), .B(n89), .C(n122), .D(\jmp_i<12> ), .Y(n191)
         );
  AOI22X1 U200 ( .A(\pc_inc_two<12> ), .B(n196), .C(\br_pre<12> ), .D(n195), 
        .Y(n190) );
  AOI22X1 U201 ( .A(n89), .B(\jmp_d<13> ), .C(n122), .D(\jmp_i<13> ), .Y(n193)
         );
  AOI22X1 U202 ( .A(\pc_inc_two<13> ), .B(n196), .C(\br_pre<13> ), .D(n195), 
        .Y(n192) );
  NAND3X1 U203 ( .A(n194), .B(n117), .C(n111), .Y(n203) );
  AOI22X1 U204 ( .A(n122), .B(\jmp_i<15> ), .C(\pc_inc_two<15> ), .D(n196), 
        .Y(n197) );
  NAND3X1 U205 ( .A(n143), .B(n145), .C(n146), .Y(n198) );
  NAND3X1 U206 ( .A(n145), .B(n143), .C(n146), .Y(\pc_nx<15> ) );
endmodule


module reg16_init ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101;

  dff_647 d0 ( .q(\read<0> ), .d(n30), .clk(clk), .rst(1'b0) );
  dff_646 d1 ( .q(\read<1> ), .d(n28), .clk(clk), .rst(1'b0) );
  dff_645 d2 ( .q(\read<2> ), .d(n26), .clk(clk), .rst(1'b0) );
  dff_644 d3 ( .q(\read<3> ), .d(n24), .clk(clk), .rst(1'b0) );
  dff_643 d4 ( .q(\read<4> ), .d(n22), .clk(clk), .rst(1'b0) );
  dff_642 d5 ( .q(\read<5> ), .d(n38), .clk(clk), .rst(1'b0) );
  dff_641 d6 ( .q(\read<6> ), .d(n20), .clk(clk), .rst(1'b0) );
  dff_640 d7 ( .q(\read<7> ), .d(n18), .clk(clk), .rst(1'b0) );
  dff_639 d8 ( .q(\read<8> ), .d(n16), .clk(clk), .rst(1'b0) );
  dff_638 d9 ( .q(\read<9> ), .d(n14), .clk(clk), .rst(1'b0) );
  dff_637 d10 ( .q(\read<10> ), .d(n12), .clk(clk), .rst(1'b0) );
  dff_636 d11 ( .q(\read<11> ), .d(n10), .clk(clk), .rst(1'b0) );
  dff_635 d12 ( .q(\read<12> ), .d(n8), .clk(clk), .rst(1'b0) );
  dff_634 d13 ( .q(\read<13> ), .d(n6), .clk(clk), .rst(1'b0) );
  dff_633 d14 ( .q(\read<14> ), .d(n4), .clk(clk), .rst(1'b0) );
  dff_632 d15 ( .q(\read<15> ), .d(n2), .clk(clk), .rst(1'b0) );
  INVX1 U3 ( .A(n98), .Y(n101) );
  OR2X1 U4 ( .A(rst), .B(wr_en), .Y(n98) );
  AND2X2 U5 ( .A(n74), .B(n46), .Y(n1) );
  INVX1 U6 ( .A(n1), .Y(n2) );
  AND2X2 U7 ( .A(n76), .B(n48), .Y(n3) );
  INVX1 U8 ( .A(n3), .Y(n4) );
  AND2X2 U9 ( .A(n78), .B(n50), .Y(n5) );
  INVX1 U10 ( .A(n5), .Y(n6) );
  AND2X2 U11 ( .A(n32), .B(n52), .Y(n7) );
  INVX1 U12 ( .A(n7), .Y(n8) );
  AND2X2 U13 ( .A(n54), .B(n41), .Y(n9) );
  INVX1 U14 ( .A(n9), .Y(n10) );
  AND2X2 U15 ( .A(n80), .B(n56), .Y(n11) );
  INVX1 U16 ( .A(n11), .Y(n12) );
  AND2X2 U17 ( .A(n34), .B(n58), .Y(n13) );
  INVX1 U18 ( .A(n13), .Y(n14) );
  AND2X2 U19 ( .A(n82), .B(n60), .Y(n15) );
  INVX1 U20 ( .A(n15), .Y(n16) );
  AND2X2 U21 ( .A(n36), .B(n62), .Y(n17) );
  INVX1 U22 ( .A(n17), .Y(n18) );
  AND2X2 U23 ( .A(n84), .B(n64), .Y(n19) );
  INVX1 U24 ( .A(n19), .Y(n20) );
  AND2X2 U25 ( .A(n88), .B(n66), .Y(n21) );
  INVX1 U26 ( .A(n21), .Y(n22) );
  AND2X2 U27 ( .A(n90), .B(n68), .Y(n23) );
  INVX1 U28 ( .A(n23), .Y(n24) );
  AND2X2 U29 ( .A(n92), .B(n70), .Y(n25) );
  INVX1 U30 ( .A(n25), .Y(n26) );
  AND2X2 U31 ( .A(n94), .B(n72), .Y(n27) );
  INVX1 U32 ( .A(n27), .Y(n28) );
  AND2X2 U33 ( .A(n96), .B(n40), .Y(n29) );
  INVX1 U34 ( .A(n29), .Y(n30) );
  AND2X2 U35 ( .A(n97), .B(\write<12> ), .Y(n31) );
  INVX1 U36 ( .A(n31), .Y(n32) );
  AND2X2 U37 ( .A(n97), .B(\write<9> ), .Y(n33) );
  INVX1 U38 ( .A(n33), .Y(n34) );
  AND2X2 U39 ( .A(n97), .B(\write<7> ), .Y(n35) );
  INVX1 U40 ( .A(n35), .Y(n36) );
  AND2X2 U41 ( .A(n86), .B(n43), .Y(n37) );
  INVX1 U42 ( .A(n37), .Y(n38) );
  AND2X2 U43 ( .A(n97), .B(\write<0> ), .Y(n39) );
  INVX1 U44 ( .A(n39), .Y(n40) );
  BUFX2 U45 ( .A(n100), .Y(n41) );
  AND2X2 U46 ( .A(n97), .B(\write<5> ), .Y(n42) );
  INVX1 U47 ( .A(n42), .Y(n43) );
  BUFX2 U48 ( .A(\write<11> ), .Y(n44) );
  AND2X1 U49 ( .A(\write<15> ), .B(n97), .Y(n45) );
  INVX1 U50 ( .A(n45), .Y(n46) );
  AND2X1 U51 ( .A(\write<14> ), .B(n97), .Y(n47) );
  INVX1 U52 ( .A(n47), .Y(n48) );
  AND2X1 U53 ( .A(\write<13> ), .B(n97), .Y(n49) );
  INVX1 U54 ( .A(n49), .Y(n50) );
  AND2X1 U55 ( .A(\read<12> ), .B(n101), .Y(n51) );
  INVX1 U56 ( .A(n51), .Y(n52) );
  AND2X1 U57 ( .A(\read<11> ), .B(n101), .Y(n53) );
  INVX1 U58 ( .A(n53), .Y(n54) );
  AND2X1 U59 ( .A(\write<10> ), .B(n97), .Y(n55) );
  INVX1 U60 ( .A(n55), .Y(n56) );
  AND2X1 U61 ( .A(\read<9> ), .B(n101), .Y(n57) );
  INVX1 U62 ( .A(n57), .Y(n58) );
  AND2X1 U63 ( .A(\write<8> ), .B(n97), .Y(n59) );
  INVX1 U64 ( .A(n59), .Y(n60) );
  AND2X1 U65 ( .A(\read<7> ), .B(n101), .Y(n61) );
  INVX1 U66 ( .A(n61), .Y(n62) );
  AND2X1 U67 ( .A(\write<6> ), .B(n97), .Y(n63) );
  INVX1 U68 ( .A(n63), .Y(n64) );
  AND2X1 U69 ( .A(\read<4> ), .B(n101), .Y(n65) );
  INVX1 U70 ( .A(n65), .Y(n66) );
  AND2X1 U71 ( .A(\write<3> ), .B(n97), .Y(n67) );
  INVX1 U72 ( .A(n67), .Y(n68) );
  AND2X1 U73 ( .A(\read<2> ), .B(n101), .Y(n69) );
  INVX1 U74 ( .A(n69), .Y(n70) );
  AND2X1 U75 ( .A(\write<1> ), .B(n97), .Y(n71) );
  INVX1 U76 ( .A(n71), .Y(n72) );
  AND2X1 U77 ( .A(\read<15> ), .B(n101), .Y(n73) );
  INVX1 U78 ( .A(n73), .Y(n74) );
  AND2X1 U79 ( .A(\read<14> ), .B(n101), .Y(n75) );
  INVX1 U80 ( .A(n75), .Y(n76) );
  AND2X1 U81 ( .A(\read<13> ), .B(n101), .Y(n77) );
  INVX1 U82 ( .A(n77), .Y(n78) );
  AND2X1 U83 ( .A(\read<10> ), .B(n101), .Y(n79) );
  INVX1 U84 ( .A(n79), .Y(n80) );
  AND2X1 U85 ( .A(\read<8> ), .B(n101), .Y(n81) );
  INVX1 U86 ( .A(n81), .Y(n82) );
  AND2X1 U87 ( .A(\read<6> ), .B(n101), .Y(n83) );
  INVX1 U88 ( .A(n83), .Y(n84) );
  AND2X1 U89 ( .A(\read<5> ), .B(n101), .Y(n85) );
  INVX1 U90 ( .A(n85), .Y(n86) );
  AND2X1 U91 ( .A(\write<4> ), .B(n97), .Y(n87) );
  INVX1 U92 ( .A(n87), .Y(n88) );
  AND2X1 U93 ( .A(\read<3> ), .B(n101), .Y(n89) );
  INVX1 U94 ( .A(n89), .Y(n90) );
  AND2X1 U95 ( .A(\write<2> ), .B(n97), .Y(n91) );
  INVX1 U96 ( .A(n91), .Y(n92) );
  AND2X1 U97 ( .A(\read<1> ), .B(n101), .Y(n93) );
  INVX1 U98 ( .A(n93), .Y(n94) );
  AND2X1 U99 ( .A(\read<0> ), .B(n101), .Y(n95) );
  INVX1 U100 ( .A(n95), .Y(n96) );
  AND2X1 U101 ( .A(wr_en), .B(n99), .Y(n97) );
  INVX1 U102 ( .A(rst), .Y(n99) );
  AOI21X1 U103 ( .A(n97), .B(n44), .C(rst), .Y(n100) );
endmodule


module reg16_35 ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54;

  dff_631 d0 ( .q(\read<0> ), .d(n39), .clk(clk), .rst(rst) );
  dff_630 d1 ( .q(\read<1> ), .d(n40), .clk(clk), .rst(rst) );
  dff_629 d2 ( .q(\read<2> ), .d(n41), .clk(clk), .rst(rst) );
  dff_628 d3 ( .q(\read<3> ), .d(n42), .clk(clk), .rst(rst) );
  dff_627 d4 ( .q(\read<4> ), .d(n43), .clk(clk), .rst(rst) );
  dff_626 d5 ( .q(\read<5> ), .d(n44), .clk(clk), .rst(rst) );
  dff_625 d6 ( .q(\read<6> ), .d(n45), .clk(clk), .rst(rst) );
  dff_624 d7 ( .q(\read<7> ), .d(n46), .clk(clk), .rst(rst) );
  dff_623 d8 ( .q(\read<8> ), .d(n47), .clk(clk), .rst(rst) );
  dff_622 d9 ( .q(\read<9> ), .d(n48), .clk(clk), .rst(rst) );
  dff_621 d10 ( .q(\read<10> ), .d(n49), .clk(clk), .rst(rst) );
  dff_620 d11 ( .q(\read<11> ), .d(n50), .clk(clk), .rst(rst) );
  dff_619 d12 ( .q(\read<12> ), .d(n51), .clk(clk), .rst(rst) );
  dff_618 d13 ( .q(\read<13> ), .d(n52), .clk(clk), .rst(rst) );
  dff_617 d14 ( .q(\read<14> ), .d(n53), .clk(clk), .rst(rst) );
  dff_616 d15 ( .q(\read<15> ), .d(n54), .clk(clk), .rst(rst) );
  INVX1 U1 ( .A(wr_en), .Y(n6) );
  INVX1 U2 ( .A(n6), .Y(n5) );
  INVX1 U3 ( .A(n5), .Y(n3) );
  INVX1 U4 ( .A(\read<6> ), .Y(n26) );
  INVX1 U5 ( .A(\read<7> ), .Y(n24) );
  INVX1 U6 ( .A(\read<10> ), .Y(n18) );
  INVX1 U7 ( .A(\read<11> ), .Y(n16) );
  INVX1 U8 ( .A(wr_en), .Y(n4) );
  INVX1 U9 ( .A(\read<12> ), .Y(n14) );
  INVX1 U10 ( .A(\read<13> ), .Y(n12) );
  INVX1 U11 ( .A(wr_en), .Y(n2) );
  INVX1 U12 ( .A(\read<14> ), .Y(n10) );
  INVX1 U13 ( .A(\read<15> ), .Y(n8) );
  INVX1 U14 ( .A(\read<0> ), .Y(n38) );
  INVX1 U15 ( .A(\read<1> ), .Y(n36) );
  INVX1 U16 ( .A(\read<2> ), .Y(n34) );
  INVX1 U17 ( .A(\read<3> ), .Y(n32) );
  INVX1 U18 ( .A(\read<4> ), .Y(n30) );
  INVX1 U19 ( .A(\read<5> ), .Y(n28) );
  INVX1 U20 ( .A(\read<8> ), .Y(n22) );
  INVX1 U21 ( .A(\read<9> ), .Y(n20) );
  INVX1 U22 ( .A(wr_en), .Y(n1) );
  MUX2X1 U23 ( .B(n7), .A(n8), .S(n1), .Y(n54) );
  MUX2X1 U24 ( .B(n23), .A(n24), .S(n1), .Y(n46) );
  MUX2X1 U25 ( .B(n9), .A(n10), .S(n2), .Y(n53) );
  MUX2X1 U26 ( .B(n15), .A(n16), .S(n4), .Y(n50) );
  INVX1 U27 ( .A(\write<0> ), .Y(n37) );
  INVX1 U28 ( .A(\write<2> ), .Y(n33) );
  INVX1 U29 ( .A(\write<1> ), .Y(n35) );
  INVX1 U30 ( .A(\write<4> ), .Y(n29) );
  INVX1 U31 ( .A(\write<8> ), .Y(n21) );
  MUX2X1 U32 ( .B(n19), .A(n20), .S(n3), .Y(n48) );
  MUX2X1 U33 ( .B(n13), .A(n14), .S(n4), .Y(n51) );
  INVX1 U34 ( .A(\write<5> ), .Y(n27) );
  INVX1 U35 ( .A(\write<3> ), .Y(n31) );
  MUX2X1 U36 ( .B(n17), .A(n18), .S(n2), .Y(n49) );
  INVX1 U37 ( .A(\write<12> ), .Y(n13) );
  INVX1 U38 ( .A(\write<6> ), .Y(n25) );
  INVX1 U39 ( .A(\write<9> ), .Y(n19) );
  MUX2X1 U40 ( .B(n11), .A(n12), .S(n1), .Y(n52) );
  INVX1 U41 ( .A(\write<10> ), .Y(n17) );
  INVX1 U42 ( .A(\write<13> ), .Y(n11) );
  INVX1 U43 ( .A(\write<7> ), .Y(n23) );
  INVX1 U44 ( .A(\write<14> ), .Y(n9) );
  INVX1 U45 ( .A(\write<15> ), .Y(n7) );
  INVX1 U46 ( .A(\write<11> ), .Y(n15) );
  MUX2X1 U47 ( .B(n22), .A(n21), .S(n5), .Y(n47) );
  MUX2X1 U48 ( .B(n26), .A(n25), .S(n5), .Y(n45) );
  MUX2X1 U49 ( .B(n28), .A(n27), .S(n5), .Y(n44) );
  MUX2X1 U50 ( .B(n30), .A(n29), .S(n5), .Y(n43) );
  MUX2X1 U51 ( .B(n32), .A(n31), .S(n5), .Y(n42) );
  MUX2X1 U52 ( .B(n34), .A(n33), .S(n5), .Y(n41) );
  MUX2X1 U53 ( .B(n36), .A(n35), .S(n5), .Y(n40) );
  MUX2X1 U54 ( .B(n38), .A(n37), .S(n5), .Y(n39) );
endmodule


module reg16_34 ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n1, n18, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86;

  dff_615 d0 ( .q(\read<0> ), .d(n86), .clk(clk), .rst(rst) );
  dff_614 d1 ( .q(\read<1> ), .d(n85), .clk(clk), .rst(rst) );
  dff_613 d2 ( .q(\read<2> ), .d(n84), .clk(clk), .rst(rst) );
  dff_612 d3 ( .q(\read<3> ), .d(n83), .clk(clk), .rst(rst) );
  dff_611 d4 ( .q(\read<4> ), .d(n82), .clk(clk), .rst(rst) );
  dff_610 d5 ( .q(\read<5> ), .d(n81), .clk(clk), .rst(rst) );
  dff_609 d6 ( .q(\read<6> ), .d(n80), .clk(clk), .rst(rst) );
  dff_608 d7 ( .q(\read<7> ), .d(n79), .clk(clk), .rst(rst) );
  dff_607 d8 ( .q(\read<8> ), .d(n78), .clk(clk), .rst(rst) );
  dff_606 d9 ( .q(\read<9> ), .d(n77), .clk(clk), .rst(rst) );
  dff_605 d10 ( .q(\read<10> ), .d(n76), .clk(clk), .rst(rst) );
  dff_604 d11 ( .q(\read<11> ), .d(n75), .clk(clk), .rst(rst) );
  dff_603 d12 ( .q(\read<12> ), .d(n74), .clk(clk), .rst(rst) );
  dff_602 d13 ( .q(\read<13> ), .d(n73), .clk(clk), .rst(rst) );
  dff_601 d14 ( .q(\read<14> ), .d(n72), .clk(clk), .rst(rst) );
  dff_600 d15 ( .q(\read<15> ), .d(n71), .clk(clk), .rst(rst) );
  AOI22X1 U18 ( .A(\read<9> ), .B(n53), .C(\write<9> ), .D(n51), .Y(n70) );
  AOI22X1 U19 ( .A(\read<8> ), .B(n53), .C(\write<8> ), .D(n51), .Y(n69) );
  AOI22X1 U20 ( .A(\read<7> ), .B(n53), .C(\write<7> ), .D(n51), .Y(n68) );
  AOI22X1 U21 ( .A(\read<6> ), .B(n53), .C(\write<6> ), .D(n51), .Y(n67) );
  AOI22X1 U22 ( .A(\read<5> ), .B(n54), .C(\write<5> ), .D(n51), .Y(n66) );
  AOI22X1 U23 ( .A(\read<4> ), .B(n54), .C(\write<4> ), .D(n51), .Y(n65) );
  AOI22X1 U24 ( .A(\read<3> ), .B(n54), .C(\write<3> ), .D(n51), .Y(n64) );
  AOI22X1 U25 ( .A(\read<2> ), .B(n54), .C(\write<2> ), .D(n51), .Y(n63) );
  AOI22X1 U26 ( .A(\read<1> ), .B(n54), .C(\write<1> ), .D(n51), .Y(n62) );
  AOI22X1 U27 ( .A(\read<15> ), .B(n54), .C(\write<15> ), .D(n51), .Y(n61) );
  AOI22X1 U28 ( .A(\read<14> ), .B(n54), .C(\write<14> ), .D(n51), .Y(n60) );
  AOI22X1 U29 ( .A(\read<13> ), .B(n54), .C(\write<13> ), .D(n51), .Y(n59) );
  AOI22X1 U30 ( .A(\read<12> ), .B(n54), .C(\write<12> ), .D(n52), .Y(n58) );
  AOI22X1 U31 ( .A(\read<11> ), .B(n54), .C(\write<11> ), .D(n52), .Y(n57) );
  AOI22X1 U32 ( .A(\read<10> ), .B(n54), .C(\write<10> ), .D(n52), .Y(n56) );
  AOI22X1 U33 ( .A(\read<0> ), .B(n54), .C(\write<0> ), .D(n52), .Y(n55) );
  INVX1 U1 ( .A(wr_en), .Y(n50) );
  INVX1 U2 ( .A(n49), .Y(n53) );
  INVX1 U3 ( .A(n50), .Y(n49) );
  INVX1 U4 ( .A(n49), .Y(n54) );
  INVX1 U5 ( .A(n53), .Y(n52) );
  INVX1 U6 ( .A(n53), .Y(n51) );
  BUFX2 U7 ( .A(n55), .Y(n1) );
  INVX1 U8 ( .A(n1), .Y(n86) );
  BUFX2 U9 ( .A(n56), .Y(n18) );
  INVX1 U10 ( .A(n18), .Y(n76) );
  BUFX2 U11 ( .A(n57), .Y(n35) );
  INVX1 U12 ( .A(n35), .Y(n75) );
  BUFX2 U13 ( .A(n58), .Y(n36) );
  INVX1 U14 ( .A(n36), .Y(n74) );
  BUFX2 U15 ( .A(n59), .Y(n37) );
  INVX1 U16 ( .A(n37), .Y(n73) );
  BUFX2 U17 ( .A(n60), .Y(n38) );
  INVX1 U34 ( .A(n38), .Y(n72) );
  BUFX2 U35 ( .A(n61), .Y(n39) );
  INVX1 U36 ( .A(n39), .Y(n71) );
  BUFX2 U37 ( .A(n62), .Y(n40) );
  INVX1 U38 ( .A(n40), .Y(n85) );
  BUFX2 U39 ( .A(n63), .Y(n41) );
  INVX1 U40 ( .A(n41), .Y(n84) );
  BUFX2 U41 ( .A(n64), .Y(n42) );
  INVX1 U42 ( .A(n42), .Y(n83) );
  BUFX2 U43 ( .A(n65), .Y(n43) );
  INVX1 U44 ( .A(n43), .Y(n82) );
  BUFX2 U45 ( .A(n66), .Y(n44) );
  INVX1 U46 ( .A(n44), .Y(n81) );
  BUFX2 U47 ( .A(n67), .Y(n45) );
  INVX1 U48 ( .A(n45), .Y(n80) );
  BUFX2 U49 ( .A(n68), .Y(n46) );
  INVX1 U50 ( .A(n46), .Y(n79) );
  BUFX2 U51 ( .A(n69), .Y(n47) );
  INVX1 U52 ( .A(n47), .Y(n78) );
  BUFX2 U53 ( .A(n70), .Y(n48) );
  INVX1 U54 ( .A(n48), .Y(n77) );
endmodule


module reg1_25 ( d, q, clk, rst, en );
  input d, clk, rst, en;
  output q;
  wire   n1, n2, n3;

  dff_599 d0 ( .q(q), .d(n3), .clk(clk), .rst(rst) );
  INVX1 U1 ( .A(q), .Y(n2) );
  INVX1 U2 ( .A(d), .Y(n1) );
  MUX2X1 U3 ( .B(n2), .A(n1), .S(en), .Y(n3) );
endmodule


module reg1_24 ( d, q, clk, rst, en );
  input d, clk, rst, en;
  output q;
  wire   n1, n2, n3;

  dff_598 d0 ( .q(q), .d(n3), .clk(clk), .rst(rst) );
  INVX1 U1 ( .A(q), .Y(n2) );
  INVX1 U2 ( .A(d), .Y(n1) );
  MUX2X1 U3 ( .B(n2), .A(n1), .S(en), .Y(n3) );
endmodule


module ID_control ( Rt_Rd, Halt, jmp_r, .opcode({\opcode<4> , \opcode<3> , 
        \opcode<2> , \opcode<1> , \opcode<0> }) );
  input \opcode<4> , \opcode<3> , \opcode<2> , \opcode<1> , \opcode<0> ;
  output Rt_Rd, Halt, jmp_r;
  wire   n3, n4, n5, n6, n7, n8, n1, n2;

  OR2X2 U3 ( .A(\opcode<2> ), .B(\opcode<3> ), .Y(n6) );
  NOR3X1 U7 ( .A(n6), .B(n3), .C(n7), .Y(Rt_Rd) );
  XOR2X1 U8 ( .A(\opcode<1> ), .B(\opcode<0> ), .Y(n7) );
  NOR3X1 U9 ( .A(n2), .B(\opcode<1> ), .C(\opcode<0> ), .Y(Halt) );
  NAND3X1 U10 ( .A(n4), .B(n3), .C(n8), .Y(n5) );
  XNOR2X1 U11 ( .A(\opcode<2> ), .B(\opcode<0> ), .Y(n8) );
  INVX1 U2 ( .A(\opcode<3> ), .Y(n4) );
  AND2X1 U4 ( .A(n1), .B(\opcode<0> ), .Y(jmp_r) );
  INVX1 U5 ( .A(\opcode<4> ), .Y(n3) );
  INVX1 U6 ( .A(n2), .Y(n1) );
  BUFX2 U12 ( .A(n5), .Y(n2) );
endmodule


module decoder ( .inst({\inst<15> , \inst<14> , \inst<13> , \inst<12> , 
        \inst<11> , \inst<10> , \inst<9> , \inst<8> , \inst<7> , \inst<6> , 
        \inst<5> , \inst<4> , \inst<3> , \inst<2> , \inst<1> , \inst<0> }), 
    .rt({\rt<2> , \rt<1> , \rt<0> }), .rs({\rs<2> , \rs<1> , \rs<0> }), .rd({
        \rd<2> , \rd<1> , \rd<0> }), .imm({\imm<15> , \imm<14> , \imm<13> , 
        \imm<12> , \imm<11> , \imm<10> , \imm<9> , \imm<8> , \imm<7> , 
        \imm<6> , \imm<5> , \imm<4> , \imm<3> , \imm<2> , \imm<1> , \imm<0> }), 
    .displacement({\displacement<15> , \displacement<14> , \displacement<13> , 
        \displacement<12> , \displacement<11> , \displacement<10> , 
        \displacement<9> , \displacement<8> , \displacement<7> , 
        \displacement<6> , \displacement<5> , \displacement<4> , 
        \displacement<3> , \displacement<2> , \displacement<1> , 
        \displacement<0> }) );
  input \inst<15> , \inst<14> , \inst<13> , \inst<12> , \inst<11> , \inst<10> ,
         \inst<9> , \inst<8> , \inst<7> , \inst<6> , \inst<5> , \inst<4> ,
         \inst<3> , \inst<2> , \inst<1> , \inst<0> ;
  output \rt<2> , \rt<1> , \rt<0> , \rs<2> , \rs<1> , \rs<0> , \rd<2> ,
         \rd<1> , \rd<0> , \imm<15> , \imm<14> , \imm<13> , \imm<12> ,
         \imm<11> , \imm<10> , \imm<9> , \imm<8> , \imm<7> , \imm<6> ,
         \imm<5> , \imm<4> , \imm<3> , \imm<2> , \imm<1> , \imm<0> ,
         \displacement<15> , \displacement<14> , \displacement<13> ,
         \displacement<12> , \displacement<11> , \displacement<10> ,
         \displacement<9> , \displacement<8> , \displacement<7> ,
         \displacement<6> , \displacement<5> , \displacement<4> ,
         \displacement<3> , \displacement<2> , \displacement<1> ,
         \displacement<0> ;
  wire   n2, n8, n9, n10, n11, n12, n14, n15, n16, n17, n20, n21, n22, n23,
         n26, n27, n28, n29, n30, n31, n34, n35, n36, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n6, n7, n13, n18, n19, n24, n25, n32, n33, n37,
         n38, n39, n49, n50, n51, n52, n53, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79;
  assign \displacement<11>  = 1'b0;
  assign \displacement<12>  = 1'b0;
  assign \displacement<13>  = 1'b0;
  assign \displacement<14>  = 1'b0;
  assign \displacement<15>  = 1'b0;

  AND2X2 U5 ( .A(n23), .B(\inst<12> ), .Y(n28) );
  NOR2X1 U39 ( .A(n15), .B(n2), .Y(\rt<2> ) );
  NOR2X1 U40 ( .A(n16), .B(n2), .Y(\rt<1> ) );
  NOR2X1 U41 ( .A(n17), .B(n2), .Y(\rt<0> ) );
  AOI21X1 U43 ( .A(n23), .B(\inst<11> ), .C(n13), .Y(n22) );
  OAI21X1 U44 ( .A(n7), .B(n15), .C(n39), .Y(\rd<2> ) );
  AOI21X1 U45 ( .A(\inst<4> ), .B(n27), .C(n28), .Y(n26) );
  OAI21X1 U46 ( .A(n7), .B(n16), .C(n38), .Y(\rd<1> ) );
  AOI21X1 U47 ( .A(\inst<3> ), .B(n27), .C(n28), .Y(n29) );
  OAI21X1 U48 ( .A(n7), .B(n17), .C(n37), .Y(\rd<0> ) );
  AOI21X1 U49 ( .A(\inst<2> ), .B(n27), .C(n28), .Y(n30) );
  OAI21X1 U50 ( .A(n14), .B(n78), .C(n2), .Y(n27) );
  OAI21X1 U51 ( .A(n78), .B(n12), .C(n60), .Y(n31) );
  NAND3X1 U52 ( .A(\inst<15> ), .B(\inst<14> ), .C(\inst<13> ), .Y(n21) );
  NAND3X1 U55 ( .A(n8), .B(\inst<7> ), .C(n73), .Y(n34) );
  OAI21X1 U56 ( .A(n69), .B(n16), .C(n71), .Y(\imm<6> ) );
  OAI21X1 U57 ( .A(n69), .B(n17), .C(n71), .Y(\imm<5> ) );
  AOI21X1 U58 ( .A(n8), .B(n73), .C(n68), .Y(n36) );
  AOI21X1 U59 ( .A(n68), .B(\inst<7> ), .C(n72), .Y(n35) );
  OAI21X1 U61 ( .A(\inst<12> ), .B(n65), .C(n33), .Y(n40) );
  AOI21X1 U62 ( .A(n8), .B(n74), .C(n62), .Y(n42) );
  NAND3X1 U68 ( .A(\inst<15> ), .B(n10), .C(\inst<13> ), .Y(n43) );
  NAND3X1 U69 ( .A(n11), .B(n9), .C(\inst<14> ), .Y(n41) );
  NAND3X1 U70 ( .A(n11), .B(n10), .C(\inst<15> ), .Y(n44) );
  NAND3X1 U71 ( .A(\inst<14> ), .B(n9), .C(\inst<13> ), .Y(n46) );
  AOI21X1 U72 ( .A(\inst<11> ), .B(n23), .C(n47), .Y(n45) );
  NOR3X1 U73 ( .A(\inst<11> ), .B(\inst<12> ), .C(n78), .Y(n47) );
  NAND3X1 U74 ( .A(\inst<14> ), .B(n11), .C(\inst<15> ), .Y(n20) );
  NOR3X1 U76 ( .A(\inst<14> ), .B(\inst<15> ), .C(n11), .Y(n23) );
  INVX1 U7 ( .A(\inst<11> ), .Y(n14) );
  AND2X1 U8 ( .A(n61), .B(n18), .Y(n75) );
  AND2X1 U9 ( .A(n23), .B(n14), .Y(n48) );
  AND2X1 U10 ( .A(n61), .B(n58), .Y(n67) );
  AND2X1 U11 ( .A(\inst<8> ), .B(n24), .Y(\rs<0> ) );
  AND2X1 U12 ( .A(\inst<9> ), .B(n24), .Y(\rs<1> ) );
  AND2X1 U13 ( .A(\inst<10> ), .B(n24), .Y(\rs<2> ) );
  AND2X1 U14 ( .A(n76), .B(\inst<0> ), .Y(\imm<0> ) );
  AND2X1 U15 ( .A(n76), .B(\inst<1> ), .Y(\imm<1> ) );
  AND2X1 U16 ( .A(n76), .B(\inst<2> ), .Y(\imm<2> ) );
  AND2X1 U17 ( .A(n76), .B(\inst<3> ), .Y(\imm<3> ) );
  AND2X1 U18 ( .A(n76), .B(\inst<4> ), .Y(\imm<4> ) );
  AND2X1 U19 ( .A(n32), .B(n64), .Y(n53) );
  AND2X1 U20 ( .A(n48), .B(\inst<0> ), .Y(\displacement<0> ) );
  AND2X1 U21 ( .A(n48), .B(\inst<1> ), .Y(\displacement<1> ) );
  AND2X1 U22 ( .A(n48), .B(\inst<2> ), .Y(\displacement<2> ) );
  AND2X1 U23 ( .A(n48), .B(\inst<3> ), .Y(\displacement<3> ) );
  AND2X1 U24 ( .A(n48), .B(\inst<4> ), .Y(\displacement<4> ) );
  AND2X1 U25 ( .A(n48), .B(\inst<5> ), .Y(\displacement<5> ) );
  AND2X1 U26 ( .A(n48), .B(\inst<6> ), .Y(\displacement<6> ) );
  AND2X1 U27 ( .A(n48), .B(\inst<7> ), .Y(\displacement<7> ) );
  AND2X1 U28 ( .A(n48), .B(\inst<8> ), .Y(\displacement<8> ) );
  AND2X1 U29 ( .A(n48), .B(\inst<9> ), .Y(\displacement<9> ) );
  AND2X1 U30 ( .A(n48), .B(\inst<10> ), .Y(\displacement<10> ) );
  INVX1 U31 ( .A(n64), .Y(\imm<8> ) );
  INVX1 U32 ( .A(\inst<5> ), .Y(n17) );
  INVX1 U33 ( .A(\inst<6> ), .Y(n16) );
  INVX1 U34 ( .A(n31), .Y(n2) );
  INVX1 U35 ( .A(\inst<12> ), .Y(n12) );
  INVX1 U36 ( .A(\inst<7> ), .Y(n15) );
  INVX1 U37 ( .A(\inst<15> ), .Y(n9) );
  INVX1 U38 ( .A(\inst<13> ), .Y(n11) );
  INVX1 U42 ( .A(\inst<14> ), .Y(n10) );
  AND2X1 U53 ( .A(n52), .B(n50), .Y(n6) );
  INVX1 U54 ( .A(n6), .Y(n7) );
  OR2X1 U60 ( .A(n66), .B(n19), .Y(n13) );
  INVX1 U63 ( .A(n13), .Y(n18) );
  OR2X1 U64 ( .A(n57), .B(n8), .Y(n19) );
  OR2X1 U65 ( .A(n77), .B(n25), .Y(n24) );
  OR2X1 U66 ( .A(n70), .B(n59), .Y(n25) );
  BUFX2 U67 ( .A(n34), .Y(n32) );
  BUFX2 U77 ( .A(n42), .Y(n33) );
  BUFX2 U78 ( .A(n30), .Y(n37) );
  BUFX2 U79 ( .A(n29), .Y(n38) );
  BUFX2 U80 ( .A(n26), .Y(n39) );
  AND2X1 U81 ( .A(n56), .B(n73), .Y(n49) );
  INVX1 U82 ( .A(n49), .Y(n50) );
  AND2X1 U83 ( .A(n56), .B(n55), .Y(n51) );
  INVX1 U84 ( .A(n51), .Y(n52) );
  INVX1 U85 ( .A(n53), .Y(\imm<7> ) );
  BUFX2 U86 ( .A(n44), .Y(n55) );
  AND2X1 U87 ( .A(n65), .B(n63), .Y(n56) );
  INVX1 U88 ( .A(n56), .Y(n57) );
  BUFX2 U89 ( .A(n46), .Y(n58) );
  INVX1 U90 ( .A(n60), .Y(n59) );
  BUFX2 U91 ( .A(n21), .Y(n60) );
  BUFX2 U92 ( .A(n45), .Y(n61) );
  INVX1 U93 ( .A(n63), .Y(n62) );
  BUFX2 U94 ( .A(n43), .Y(n63) );
  BUFX2 U95 ( .A(n35), .Y(n64) );
  BUFX2 U96 ( .A(n41), .Y(n65) );
  INVX1 U97 ( .A(n58), .Y(n66) );
  INVX1 U98 ( .A(n67), .Y(n68) );
  BUFX2 U99 ( .A(n36), .Y(n69) );
  INVX1 U100 ( .A(n22), .Y(n70) );
  INVX1 U101 ( .A(n72), .Y(n71) );
  AND2X1 U102 ( .A(\inst<4> ), .B(n40), .Y(n72) );
  AND2X1 U103 ( .A(\inst<12> ), .B(n14), .Y(n73) );
  INVX1 U104 ( .A(n73), .Y(n74) );
  INVX1 U105 ( .A(n55), .Y(n8) );
  INVX1 U106 ( .A(n75), .Y(n76) );
  INVX1 U107 ( .A(n78), .Y(n77) );
  BUFX2 U108 ( .A(n20), .Y(n78) );
  INVX1 U109 ( .A(n79), .Y(\imm<9> ) );
  INVX1 U110 ( .A(n79), .Y(\imm<10> ) );
  INVX1 U111 ( .A(n79), .Y(\imm<11> ) );
  INVX1 U112 ( .A(n79), .Y(\imm<12> ) );
  INVX1 U113 ( .A(n79), .Y(\imm<13> ) );
  INVX1 U114 ( .A(n79), .Y(\imm<14> ) );
  INVX1 U115 ( .A(n79), .Y(\imm<15> ) );
  INVX1 U116 ( .A(\imm<8> ), .Y(n79) );
endmodule


module rf_bypass ( .read1data({\read1data<15> , \read1data<14> , 
        \read1data<13> , \read1data<12> , \read1data<11> , \read1data<10> , 
        \read1data<9> , \read1data<8> , \read1data<7> , \read1data<6> , 
        \read1data<5> , \read1data<4> , \read1data<3> , \read1data<2> , 
        \read1data<1> , \read1data<0> }), .read2data({\read2data<15> , 
        \read2data<14> , \read2data<13> , \read2data<12> , \read2data<11> , 
        \read2data<10> , \read2data<9> , \read2data<8> , \read2data<7> , 
        \read2data<6> , \read2data<5> , \read2data<4> , \read2data<3> , 
        \read2data<2> , \read2data<1> , \read2data<0> }), err, clk, rst, 
    .read1regsel({\read1regsel<2> , \read1regsel<1> , \read1regsel<0> }), 
    .read2regsel({\read2regsel<2> , \read2regsel<1> , \read2regsel<0> }), 
    .writeregsel({\writeregsel<2> , \writeregsel<1> , \writeregsel<0> }), 
    .writedata({\writedata<15> , \writedata<14> , \writedata<13> , 
        \writedata<12> , \writedata<11> , \writedata<10> , \writedata<9> , 
        \writedata<8> , \writedata<7> , \writedata<6> , \writedata<5> , 
        \writedata<4> , \writedata<3> , \writedata<2> , \writedata<1> , 
        \writedata<0> }), write );
  input clk, rst, \read1regsel<2> , \read1regsel<1> , \read1regsel<0> ,
         \read2regsel<2> , \read2regsel<1> , \read2regsel<0> ,
         \writeregsel<2> , \writeregsel<1> , \writeregsel<0> , \writedata<15> ,
         \writedata<14> , \writedata<13> , \writedata<12> , \writedata<11> ,
         \writedata<10> , \writedata<9> , \writedata<8> , \writedata<7> ,
         \writedata<6> , \writedata<5> , \writedata<4> , \writedata<3> ,
         \writedata<2> , \writedata<1> , \writedata<0> , write;
  output \read1data<15> , \read1data<14> , \read1data<13> , \read1data<12> ,
         \read1data<11> , \read1data<10> , \read1data<9> , \read1data<8> ,
         \read1data<7> , \read1data<6> , \read1data<5> , \read1data<4> ,
         \read1data<3> , \read1data<2> , \read1data<1> , \read1data<0> ,
         \read2data<15> , \read2data<14> , \read2data<13> , \read2data<12> ,
         \read2data<11> , \read2data<10> , \read2data<9> , \read2data<8> ,
         \read2data<7> , \read2data<6> , \read2data<5> , \read2data<4> ,
         \read2data<3> , \read2data<2> , \read2data<1> , \read2data<0> , err;
  wire   n109, \read1tmp<15> , \read1tmp<14> , \read1tmp<13> , \read1tmp<12> ,
         \read1tmp<11> , \read1tmp<10> , \read1tmp<9> , \read1tmp<8> ,
         \read1tmp<7> , \read1tmp<6> , \read1tmp<5> , \read1tmp<4> ,
         \read1tmp<3> , \read1tmp<2> , \read1tmp<1> , \read1tmp<0> ,
         \read2tmp<15> , \read2tmp<14> , \read2tmp<13> , \read2tmp<12> ,
         \read2tmp<11> , \read2tmp<10> , \read2tmp<9> , \read2tmp<8> ,
         \read2tmp<7> , \read2tmp<6> , \read2tmp<5> , \read2tmp<4> ,
         \read2tmp<3> , \read2tmp<2> , \read2tmp<1> , \read2tmp<0> , n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n40, n41, n43, n44, n61, n62, n64, n1, n2, n3, n4, n5, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n42, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n63, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n103, n104, n105, n106, n107, n108;
  assign err = 1'b0;

  rf RFile ( .read1data({\read1tmp<15> , \read1tmp<14> , \read1tmp<13> , 
        \read1tmp<12> , \read1tmp<11> , \read1tmp<10> , \read1tmp<9> , 
        \read1tmp<8> , \read1tmp<7> , \read1tmp<6> , \read1tmp<5> , 
        \read1tmp<4> , \read1tmp<3> , \read1tmp<2> , \read1tmp<1> , 
        \read1tmp<0> }), .read2data({\read2tmp<15> , \read2tmp<14> , 
        \read2tmp<13> , \read2tmp<12> , \read2tmp<11> , \read2tmp<10> , 
        \read2tmp<9> , \read2tmp<8> , \read2tmp<7> , \read2tmp<6> , 
        \read2tmp<5> , \read2tmp<4> , \read2tmp<3> , \read2tmp<2> , 
        \read2tmp<1> , \read2tmp<0> }), .err(n109), .clk(clk), .rst(rst), 
        .read1regsel({\read1regsel<2> , \read1regsel<1> , \read1regsel<0> }), 
        .read2regsel({\read2regsel<2> , \read2regsel<1> , \read2regsel<0> }), 
        .writeregsel({\writeregsel<2> , \writeregsel<1> , \writeregsel<0> }), 
        .writedata({\writedata<15> , \writedata<14> , \writedata<13> , 
        \writedata<12> , \writedata<11> , \writedata<10> , \writedata<9> , 
        \writedata<8> , \writedata<7> , \writedata<6> , \writedata<5> , 
        \writedata<4> , \writedata<3> , \writedata<2> , \writedata<1> , 
        \writedata<0> }), .write(write) );
  OAI21X1 U18 ( .A(n106), .B(n12), .C(n95), .Y(\read2data<9> ) );
  OAI21X1 U20 ( .A(n106), .B(n13), .C(n93), .Y(\read2data<8> ) );
  OAI21X1 U22 ( .A(n106), .B(n14), .C(n91), .Y(\read2data<7> ) );
  OAI21X1 U24 ( .A(n106), .B(n15), .C(n89), .Y(\read2data<6> ) );
  OAI21X1 U26 ( .A(n106), .B(n16), .C(n87), .Y(\read2data<5> ) );
  OAI21X1 U28 ( .A(n106), .B(n17), .C(n85), .Y(\read2data<4> ) );
  OAI21X1 U30 ( .A(n106), .B(n18), .C(n83), .Y(\read2data<3> ) );
  OAI21X1 U32 ( .A(n106), .B(n19), .C(n81), .Y(\read2data<2> ) );
  OAI21X1 U34 ( .A(n106), .B(n20), .C(n79), .Y(\read2data<1> ) );
  OAI21X1 U36 ( .A(n106), .B(n6), .C(n77), .Y(\read2data<15> ) );
  OAI21X1 U38 ( .A(n106), .B(n7), .C(n75), .Y(\read2data<14> ) );
  OAI21X1 U40 ( .A(n106), .B(n8), .C(n73), .Y(\read2data<13> ) );
  OAI21X1 U42 ( .A(n107), .B(n9), .C(n71), .Y(\read2data<12> ) );
  OAI21X1 U44 ( .A(n107), .B(n10), .C(n67), .Y(\read2data<11> ) );
  OAI21X1 U46 ( .A(n107), .B(n11), .C(n60), .Y(\read2data<10> ) );
  OAI21X1 U48 ( .A(n107), .B(n21), .C(n56), .Y(\read2data<0> ) );
  NAND3X1 U50 ( .A(n40), .B(n41), .C(n99), .Y(n23) );
  XOR2X1 U52 ( .A(\writeregsel<2> ), .B(\read2regsel<2> ), .Y(n43) );
  XNOR2X1 U53 ( .A(\writeregsel<1> ), .B(\read2regsel<1> ), .Y(n41) );
  XNOR2X1 U54 ( .A(\writeregsel<0> ), .B(\read2regsel<0> ), .Y(n40) );
  OAI21X1 U55 ( .A(n12), .B(n103), .C(n54), .Y(\read1data<9> ) );
  OAI21X1 U57 ( .A(n13), .B(n103), .C(n52), .Y(\read1data<8> ) );
  OAI21X1 U59 ( .A(n14), .B(n103), .C(n50), .Y(\read1data<7> ) );
  OAI21X1 U61 ( .A(n15), .B(n103), .C(n48), .Y(\read1data<6> ) );
  OAI21X1 U63 ( .A(n16), .B(n103), .C(n46), .Y(\read1data<5> ) );
  OAI21X1 U65 ( .A(n17), .B(n103), .C(n42), .Y(\read1data<4> ) );
  OAI21X1 U67 ( .A(n18), .B(n103), .C(n38), .Y(\read1data<3> ) );
  OAI21X1 U69 ( .A(n19), .B(n103), .C(n36), .Y(\read1data<2> ) );
  OAI21X1 U71 ( .A(n20), .B(n103), .C(n34), .Y(\read1data<1> ) );
  OAI21X1 U73 ( .A(n6), .B(n103), .C(n32), .Y(\read1data<15> ) );
  OAI21X1 U75 ( .A(n7), .B(n103), .C(n30), .Y(\read1data<14> ) );
  OAI21X1 U77 ( .A(n8), .B(n103), .C(n28), .Y(\read1data<13> ) );
  OAI21X1 U79 ( .A(n9), .B(n104), .C(n26), .Y(\read1data<12> ) );
  OAI21X1 U81 ( .A(n10), .B(n104), .C(n24), .Y(\read1data<11> ) );
  OAI21X1 U83 ( .A(n11), .B(n104), .C(n4), .Y(\read1data<10> ) );
  OAI21X1 U85 ( .A(n21), .B(n104), .C(n2), .Y(\read1data<0> ) );
  NAND3X1 U87 ( .A(n61), .B(n62), .C(n97), .Y(n44) );
  XOR2X1 U89 ( .A(\writeregsel<2> ), .B(\read1regsel<2> ), .Y(n64) );
  XNOR2X1 U90 ( .A(\writeregsel<1> ), .B(\read1regsel<1> ), .Y(n62) );
  XNOR2X1 U91 ( .A(\writeregsel<0> ), .B(\read1regsel<0> ), .Y(n61) );
  INVX1 U1 ( .A(write), .Y(n22) );
  INVX1 U2 ( .A(\writedata<3> ), .Y(n18) );
  INVX1 U3 ( .A(\writedata<5> ), .Y(n16) );
  INVX1 U4 ( .A(\writedata<6> ), .Y(n15) );
  INVX1 U5 ( .A(\writedata<9> ), .Y(n12) );
  INVX1 U6 ( .A(\writedata<14> ), .Y(n7) );
  INVX2 U7 ( .A(n105), .Y(n103) );
  INVX2 U8 ( .A(n105), .Y(n104) );
  AND2X1 U9 ( .A(\read1tmp<0> ), .B(n104), .Y(n1) );
  INVX1 U10 ( .A(n1), .Y(n2) );
  AND2X1 U11 ( .A(\read1tmp<10> ), .B(n103), .Y(n3) );
  INVX1 U12 ( .A(n3), .Y(n4) );
  AND2X1 U13 ( .A(\read1tmp<11> ), .B(n104), .Y(n5) );
  INVX1 U14 ( .A(n5), .Y(n24) );
  AND2X1 U15 ( .A(\read1tmp<12> ), .B(n104), .Y(n25) );
  INVX1 U16 ( .A(n25), .Y(n26) );
  AND2X1 U17 ( .A(\read1tmp<13> ), .B(n104), .Y(n27) );
  INVX1 U19 ( .A(n27), .Y(n28) );
  AND2X1 U21 ( .A(\read1tmp<14> ), .B(n104), .Y(n29) );
  INVX1 U23 ( .A(n29), .Y(n30) );
  AND2X1 U25 ( .A(\read1tmp<15> ), .B(n104), .Y(n31) );
  INVX1 U27 ( .A(n31), .Y(n32) );
  AND2X1 U29 ( .A(\read1tmp<1> ), .B(n104), .Y(n33) );
  INVX1 U31 ( .A(n33), .Y(n34) );
  AND2X1 U33 ( .A(\read1tmp<2> ), .B(n104), .Y(n35) );
  INVX1 U35 ( .A(n35), .Y(n36) );
  AND2X1 U37 ( .A(\read1tmp<3> ), .B(n104), .Y(n37) );
  INVX1 U39 ( .A(n37), .Y(n38) );
  AND2X1 U41 ( .A(\read1tmp<4> ), .B(n104), .Y(n39) );
  INVX1 U43 ( .A(n39), .Y(n42) );
  AND2X1 U45 ( .A(\read1tmp<5> ), .B(n104), .Y(n45) );
  INVX1 U47 ( .A(n45), .Y(n46) );
  AND2X1 U49 ( .A(\read1tmp<6> ), .B(n104), .Y(n47) );
  INVX1 U51 ( .A(n47), .Y(n48) );
  AND2X1 U56 ( .A(\read1tmp<7> ), .B(n104), .Y(n49) );
  INVX1 U58 ( .A(n49), .Y(n50) );
  AND2X1 U60 ( .A(\read1tmp<8> ), .B(n103), .Y(n51) );
  INVX1 U62 ( .A(n51), .Y(n52) );
  AND2X1 U64 ( .A(\read1tmp<9> ), .B(n103), .Y(n53) );
  INVX1 U66 ( .A(n53), .Y(n54) );
  INVX1 U68 ( .A(n58), .Y(n55) );
  INVX1 U70 ( .A(n55), .Y(n56) );
  AND2X1 U72 ( .A(\read2tmp<0> ), .B(n106), .Y(n57) );
  INVX1 U74 ( .A(n57), .Y(n58) );
  INVX1 U76 ( .A(n65), .Y(n59) );
  INVX1 U78 ( .A(n59), .Y(n60) );
  AND2X1 U80 ( .A(\read2tmp<10> ), .B(n106), .Y(n63) );
  INVX1 U82 ( .A(n63), .Y(n65) );
  INVX1 U84 ( .A(n69), .Y(n66) );
  INVX1 U86 ( .A(n66), .Y(n67) );
  AND2X1 U88 ( .A(\read2tmp<11> ), .B(n107), .Y(n68) );
  INVX1 U92 ( .A(n68), .Y(n69) );
  AND2X1 U93 ( .A(\read2tmp<12> ), .B(n107), .Y(n70) );
  INVX1 U94 ( .A(n70), .Y(n71) );
  AND2X1 U95 ( .A(\read2tmp<13> ), .B(n107), .Y(n72) );
  INVX1 U96 ( .A(n72), .Y(n73) );
  AND2X1 U97 ( .A(\read2tmp<14> ), .B(n107), .Y(n74) );
  INVX1 U98 ( .A(n74), .Y(n75) );
  AND2X1 U99 ( .A(\read2tmp<15> ), .B(n107), .Y(n76) );
  INVX1 U100 ( .A(n76), .Y(n77) );
  AND2X1 U101 ( .A(\read2tmp<1> ), .B(n107), .Y(n78) );
  INVX1 U102 ( .A(n78), .Y(n79) );
  AND2X1 U103 ( .A(\read2tmp<2> ), .B(n107), .Y(n80) );
  INVX1 U104 ( .A(n80), .Y(n81) );
  AND2X1 U105 ( .A(\read2tmp<3> ), .B(n107), .Y(n82) );
  INVX1 U106 ( .A(n82), .Y(n83) );
  AND2X1 U107 ( .A(\read2tmp<4> ), .B(n107), .Y(n84) );
  INVX1 U108 ( .A(n84), .Y(n85) );
  AND2X1 U109 ( .A(\read2tmp<5> ), .B(n107), .Y(n86) );
  INVX1 U110 ( .A(n86), .Y(n87) );
  AND2X1 U111 ( .A(\read2tmp<6> ), .B(n107), .Y(n88) );
  INVX1 U112 ( .A(n88), .Y(n89) );
  AND2X1 U113 ( .A(\read2tmp<7> ), .B(n106), .Y(n90) );
  INVX1 U114 ( .A(n90), .Y(n91) );
  AND2X1 U115 ( .A(\read2tmp<8> ), .B(n106), .Y(n92) );
  INVX1 U116 ( .A(n92), .Y(n93) );
  AND2X1 U117 ( .A(\read2tmp<9> ), .B(n107), .Y(n94) );
  INVX1 U118 ( .A(n94), .Y(n95) );
  OR2X1 U119 ( .A(n22), .B(n64), .Y(n96) );
  INVX1 U120 ( .A(n96), .Y(n97) );
  OR2X1 U121 ( .A(n22), .B(n43), .Y(n98) );
  INVX1 U122 ( .A(n98), .Y(n99) );
  BUFX2 U123 ( .A(n44), .Y(n100) );
  INVX1 U124 ( .A(n100), .Y(n105) );
  BUFX2 U125 ( .A(n23), .Y(n101) );
  INVX1 U126 ( .A(n101), .Y(n108) );
  INVX1 U128 ( .A(\writedata<12> ), .Y(n9) );
  INVX1 U129 ( .A(\writedata<11> ), .Y(n10) );
  INVX1 U130 ( .A(\writedata<2> ), .Y(n19) );
  INVX1 U131 ( .A(\writedata<13> ), .Y(n8) );
  INVX1 U132 ( .A(\writedata<8> ), .Y(n13) );
  INVX1 U133 ( .A(\writedata<15> ), .Y(n6) );
  INVX1 U134 ( .A(\writedata<1> ), .Y(n20) );
  INVX1 U135 ( .A(\writedata<0> ), .Y(n21) );
  INVX1 U136 ( .A(\writedata<10> ), .Y(n11) );
  INVX1 U137 ( .A(\writedata<4> ), .Y(n17) );
  INVX1 U138 ( .A(\writedata<7> ), .Y(n14) );
  INVX8 U139 ( .A(n108), .Y(n106) );
  INVX8 U140 ( .A(n108), .Y(n107) );
endmodule


module reg_control ( rs_v, rt_v, rd_v, .r1_reg({\r1_reg<2> , \r1_reg<1> , 
        \r1_reg<0> }), .r2_reg({\r2_reg<2> , \r2_reg<1> , \r2_reg<0> }), 
    .r_wr({\r_wr<2> , \r_wr<1> , \r_wr<0> }), .inst({\inst<15> , \inst<14> , 
        \inst<13> , \inst<12> , \inst<11> , \inst<10> , \inst<9> , \inst<8> , 
        \inst<7> , \inst<6> , \inst<5> , \inst<4> , \inst<3> , \inst<2> , 
        \inst<1> , \inst<0> }) );
  input \inst<15> , \inst<14> , \inst<13> , \inst<12> , \inst<11> , \inst<10> ,
         \inst<9> , \inst<8> , \inst<7> , \inst<6> , \inst<5> , \inst<4> ,
         \inst<3> , \inst<2> , \inst<1> , \inst<0> ;
  output rs_v, rt_v, rd_v, \r1_reg<2> , \r1_reg<1> , \r1_reg<0> , \r2_reg<2> ,
         \r2_reg<1> , \r2_reg<0> , \r_wr<2> , \r_wr<1> , \r_wr<0> ;
  wire   n66, n67, n68, n69, n2, n3, n4, n7, n8, n9, n10, n12, n13, n14, n15,
         n17, n18, n21, n23, n24, n26, n27, n28, n29, n31, n33, n34, n36, n37,
         n1, n5, n6, n11, n16, n19, n20, n22, n25, n30, n32, n35, n38, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65;

  AND2X2 U5 ( .A(rt_v), .B(\inst<6> ), .Y(\r2_reg<1> ) );
  AND2X2 U6 ( .A(rt_v), .B(\inst<5> ), .Y(\r2_reg<0> ) );
  AND2X2 U7 ( .A(rs_v), .B(\inst<10> ), .Y(\r1_reg<2> ) );
  AND2X2 U8 ( .A(rs_v), .B(\inst<9> ), .Y(\r1_reg<1> ) );
  AND2X2 U9 ( .A(rs_v), .B(\inst<8> ), .Y(\r1_reg<0> ) );
  INVX2 U18 ( .A(\inst<11> ), .Y(n10) );
  NAND3X1 U19 ( .A(n52), .B(n64), .C(n48), .Y(n66) );
  AOI21X1 U20 ( .A(n43), .B(\inst<12> ), .C(n14), .Y(n12) );
  AOI21X1 U21 ( .A(n8), .B(n3), .C(\inst<14> ), .Y(n13) );
  NAND3X1 U22 ( .A(n35), .B(n61), .C(n47), .Y(n67) );
  AOI22X1 U23 ( .A(\inst<10> ), .B(n56), .C(\inst<7> ), .D(n2), .Y(n18) );
  NAND3X1 U25 ( .A(n30), .B(n61), .C(n46), .Y(n68) );
  AOI22X1 U26 ( .A(\inst<9> ), .B(n56), .C(\inst<6> ), .D(n2), .Y(n21) );
  NAND3X1 U28 ( .A(n22), .B(n61), .C(n45), .Y(n69) );
  AOI22X1 U29 ( .A(\inst<8> ), .B(n56), .C(\inst<5> ), .D(n2), .Y(n23) );
  AOI21X1 U30 ( .A(n4), .B(\inst<13> ), .C(n14), .Y(n24) );
  OAI21X1 U31 ( .A(n63), .B(n26), .C(n19), .Y(n14) );
  NAND3X1 U32 ( .A(n8), .B(n3), .C(\inst<14> ), .Y(n27) );
  OAI21X1 U33 ( .A(\inst<13> ), .B(\inst<11> ), .C(n9), .Y(n26) );
  NAND3X1 U36 ( .A(n4), .B(n8), .C(\inst<12> ), .Y(n28) );
  NAND3X1 U37 ( .A(\inst<13> ), .B(\inst<12> ), .C(n31), .Y(n17) );
  AOI21X1 U39 ( .A(n10), .B(n58), .C(n53), .Y(n15) );
  OAI21X1 U40 ( .A(n58), .B(n53), .C(n16), .Y(rt_v) );
  AOI21X1 U41 ( .A(n29), .B(n4), .C(n34), .Y(n33) );
  NOR3X1 U42 ( .A(n50), .B(\inst<13> ), .C(n63), .Y(n34) );
  NOR3X1 U45 ( .A(\inst<12> ), .B(\inst<13> ), .C(\inst<11> ), .Y(n29) );
  OAI21X1 U47 ( .A(\inst<15> ), .B(n7), .C(n5), .Y(rs_v) );
  AOI22X1 U48 ( .A(\inst<13> ), .B(\inst<11> ), .C(\inst<15> ), .D(n44), .Y(
        n36) );
  NAND3X1 U49 ( .A(\inst<14> ), .B(n10), .C(n58), .Y(n37) );
  INVX1 U3 ( .A(\inst<14> ), .Y(n7) );
  AND2X1 U4 ( .A(n6), .B(n52), .Y(n55) );
  INVX1 U10 ( .A(\inst<12> ), .Y(n9) );
  INVX1 U11 ( .A(\inst<15> ), .Y(n3) );
  AND2X1 U12 ( .A(rt_v), .B(\inst<7> ), .Y(\r2_reg<2> ) );
  INVX1 U13 ( .A(n36), .Y(n1) );
  INVX1 U14 ( .A(n1), .Y(n5) );
  AND2X1 U15 ( .A(n3), .B(n7), .Y(n31) );
  INVX1 U16 ( .A(\inst<13> ), .Y(n8) );
  INVX1 U17 ( .A(n63), .Y(n4) );
  BUFX2 U24 ( .A(n28), .Y(n6) );
  INVX1 U27 ( .A(n33), .Y(n11) );
  INVX1 U34 ( .A(n11), .Y(n16) );
  BUFX2 U35 ( .A(n27), .Y(n19) );
  AND2X1 U38 ( .A(\inst<2> ), .B(n65), .Y(n20) );
  INVX1 U43 ( .A(n20), .Y(n22) );
  AND2X1 U44 ( .A(\inst<3> ), .B(n65), .Y(n25) );
  INVX1 U46 ( .A(n25), .Y(n30) );
  AND2X1 U50 ( .A(\inst<4> ), .B(n65), .Y(n32) );
  INVX1 U51 ( .A(n32), .Y(n35) );
  BUFX2 U52 ( .A(n24), .Y(n38) );
  INVX1 U53 ( .A(n38), .Y(n2) );
  BUFX2 U54 ( .A(n69), .Y(\r_wr<0> ) );
  BUFX2 U55 ( .A(n68), .Y(\r_wr<1> ) );
  BUFX2 U56 ( .A(n67), .Y(\r_wr<2> ) );
  BUFX2 U57 ( .A(n66), .Y(rd_v) );
  BUFX2 U58 ( .A(n13), .Y(n43) );
  BUFX2 U59 ( .A(n37), .Y(n44) );
  BUFX2 U60 ( .A(n23), .Y(n45) );
  BUFX2 U61 ( .A(n21), .Y(n46) );
  BUFX2 U62 ( .A(n18), .Y(n47) );
  BUFX2 U63 ( .A(n12), .Y(n48) );
  AND2X1 U64 ( .A(\inst<12> ), .B(\inst<11> ), .Y(n49) );
  INVX1 U65 ( .A(n49), .Y(n50) );
  AND2X1 U66 ( .A(n54), .B(n29), .Y(n51) );
  INVX1 U67 ( .A(n51), .Y(n52) );
  INVX1 U68 ( .A(n54), .Y(n53) );
  AND2X1 U69 ( .A(\inst<14> ), .B(\inst<15> ), .Y(n54) );
  INVX1 U70 ( .A(n55), .Y(n56) );
  INVX1 U71 ( .A(n60), .Y(n57) );
  INVX1 U72 ( .A(n57), .Y(n58) );
  OR2X1 U73 ( .A(\inst<13> ), .B(\inst<12> ), .Y(n59) );
  INVX1 U74 ( .A(n59), .Y(n60) );
  BUFX2 U75 ( .A(n17), .Y(n61) );
  AND2X1 U76 ( .A(\inst<15> ), .B(n7), .Y(n62) );
  INVX1 U77 ( .A(n62), .Y(n63) );
  INVX1 U78 ( .A(n65), .Y(n64) );
  BUFX2 U79 ( .A(n15), .Y(n65) );
endmodule


module reg3_8 ( .read({\read<2> , \read<1> , \read<0> }), .write({\write<2> , 
        \write<1> , \write<0> }), wr_en, rst, clk );
  input \write<2> , \write<1> , \write<0> , wr_en, rst, clk;
  output \read<2> , \read<1> , \read<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;

  dff_597 d0 ( .q(\read<0> ), .d(n7), .clk(clk), .rst(rst) );
  dff_596 d1 ( .q(\read<1> ), .d(n8), .clk(clk), .rst(rst) );
  dff_595 d2 ( .q(\read<2> ), .d(n9), .clk(clk), .rst(rst) );
  INVX1 U1 ( .A(\read<0> ), .Y(n6) );
  INVX1 U2 ( .A(\read<1> ), .Y(n4) );
  INVX1 U3 ( .A(\read<2> ), .Y(n2) );
  INVX1 U4 ( .A(\write<0> ), .Y(n5) );
  INVX1 U5 ( .A(\write<1> ), .Y(n3) );
  INVX1 U6 ( .A(\write<2> ), .Y(n1) );
  MUX2X1 U7 ( .B(n2), .A(n1), .S(wr_en), .Y(n9) );
  MUX2X1 U8 ( .B(n4), .A(n3), .S(wr_en), .Y(n8) );
  MUX2X1 U9 ( .B(n6), .A(n5), .S(wr_en), .Y(n7) );
endmodule


module reg3_7 ( .read({\read<2> , \read<1> , \read<0> }), .write({\write<2> , 
        \write<1> , \write<0> }), wr_en, rst, clk );
  input \write<2> , \write<1> , \write<0> , wr_en, rst, clk;
  output \read<2> , \read<1> , \read<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;

  dff_594 d0 ( .q(\read<0> ), .d(n7), .clk(clk), .rst(rst) );
  dff_593 d1 ( .q(\read<1> ), .d(n8), .clk(clk), .rst(rst) );
  dff_592 d2 ( .q(\read<2> ), .d(n9), .clk(clk), .rst(rst) );
  INVX1 U1 ( .A(\read<0> ), .Y(n6) );
  INVX1 U2 ( .A(\read<1> ), .Y(n4) );
  INVX1 U3 ( .A(\read<2> ), .Y(n2) );
  INVX1 U4 ( .A(\write<0> ), .Y(n5) );
  INVX1 U5 ( .A(\write<1> ), .Y(n3) );
  INVX1 U6 ( .A(\write<2> ), .Y(n1) );
  MUX2X1 U7 ( .B(n2), .A(n1), .S(wr_en), .Y(n9) );
  MUX2X1 U8 ( .B(n4), .A(n3), .S(wr_en), .Y(n8) );
  MUX2X1 U9 ( .B(n6), .A(n5), .S(wr_en), .Y(n7) );
endmodule


module reg3_6 ( .read({\read<2> , \read<1> , \read<0> }), .write({\write<2> , 
        \write<1> , \write<0> }), wr_en, rst, clk );
  input \write<2> , \write<1> , \write<0> , wr_en, rst, clk;
  output \read<2> , \read<1> , \read<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;

  dff_591 d0 ( .q(\read<0> ), .d(n7), .clk(clk), .rst(rst) );
  dff_590 d1 ( .q(\read<1> ), .d(n8), .clk(clk), .rst(rst) );
  dff_589 d2 ( .q(\read<2> ), .d(n9), .clk(clk), .rst(rst) );
  INVX1 U1 ( .A(\read<0> ), .Y(n6) );
  INVX1 U2 ( .A(\read<1> ), .Y(n4) );
  INVX1 U3 ( .A(\read<2> ), .Y(n2) );
  INVX1 U4 ( .A(\write<0> ), .Y(n5) );
  INVX1 U5 ( .A(\write<1> ), .Y(n3) );
  INVX1 U6 ( .A(\write<2> ), .Y(n1) );
  MUX2X1 U7 ( .B(n2), .A(n1), .S(wr_en), .Y(n9) );
  MUX2X1 U8 ( .B(n4), .A(n3), .S(wr_en), .Y(n8) );
  MUX2X1 U9 ( .B(n6), .A(n5), .S(wr_en), .Y(n7) );
endmodule


module reg16_33 ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n58, n1, n2, n3, n4, n5, n6, n7, n8, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57;

  dff_588 d0 ( .q(\read<0> ), .d(n42), .clk(clk), .rst(rst) );
  dff_587 d1 ( .q(\read<1> ), .d(n43), .clk(clk), .rst(rst) );
  dff_586 d2 ( .q(\read<2> ), .d(n44), .clk(clk), .rst(rst) );
  dff_585 d3 ( .q(\read<3> ), .d(n45), .clk(clk), .rst(rst) );
  dff_584 d4 ( .q(\read<4> ), .d(n46), .clk(clk), .rst(rst) );
  dff_583 d5 ( .q(\read<5> ), .d(n47), .clk(clk), .rst(rst) );
  dff_582 d6 ( .q(\read<6> ), .d(n48), .clk(clk), .rst(rst) );
  dff_581 d7 ( .q(n58), .d(n49), .clk(clk), .rst(rst) );
  dff_580 d8 ( .q(\read<8> ), .d(n50), .clk(clk), .rst(rst) );
  dff_579 d9 ( .q(\read<9> ), .d(n51), .clk(clk), .rst(rst) );
  dff_578 d10 ( .q(\read<10> ), .d(n52), .clk(clk), .rst(rst) );
  dff_577 d11 ( .q(\read<11> ), .d(n53), .clk(clk), .rst(rst) );
  dff_576 d12 ( .q(\read<12> ), .d(n54), .clk(clk), .rst(rst) );
  dff_575 d13 ( .q(\read<13> ), .d(n55), .clk(clk), .rst(rst) );
  dff_574 d14 ( .q(\read<14> ), .d(n56), .clk(clk), .rst(rst) );
  dff_573 d15 ( .q(\read<15> ), .d(n57), .clk(clk), .rst(rst) );
  INVX1 U1 ( .A(wr_en), .Y(n8) );
  INVX1 U2 ( .A(n58), .Y(n10) );
  INVX1 U3 ( .A(n8), .Y(n6) );
  INVX1 U4 ( .A(n10), .Y(\read<7> ) );
  INVX1 U5 ( .A(n8), .Y(n7) );
  INVX1 U6 ( .A(\read<0> ), .Y(n41) );
  INVX1 U7 ( .A(\read<1> ), .Y(n39) );
  INVX1 U8 ( .A(\read<2> ), .Y(n37) );
  INVX1 U9 ( .A(\read<3> ), .Y(n35) );
  INVX1 U10 ( .A(\read<4> ), .Y(n33) );
  INVX1 U11 ( .A(\read<5> ), .Y(n31) );
  INVX1 U12 ( .A(\read<6> ), .Y(n29) );
  INVX1 U13 ( .A(\read<8> ), .Y(n26) );
  INVX1 U14 ( .A(\read<9> ), .Y(n24) );
  INVX1 U15 ( .A(\read<10> ), .Y(n22) );
  BUFX2 U16 ( .A(\read<13> ), .Y(n1) );
  BUFX2 U17 ( .A(\read<11> ), .Y(n2) );
  BUFX2 U18 ( .A(\read<14> ), .Y(n3) );
  BUFX2 U19 ( .A(\read<15> ), .Y(n4) );
  INVX1 U20 ( .A(n1), .Y(n16) );
  INVX1 U21 ( .A(n2), .Y(n20) );
  INVX1 U22 ( .A(\write<0> ), .Y(n40) );
  INVX1 U23 ( .A(\write<1> ), .Y(n38) );
  INVX1 U24 ( .A(\write<2> ), .Y(n36) );
  INVX1 U25 ( .A(\write<3> ), .Y(n34) );
  INVX1 U26 ( .A(\write<4> ), .Y(n32) );
  INVX1 U27 ( .A(\write<5> ), .Y(n30) );
  INVX1 U28 ( .A(\write<6> ), .Y(n28) );
  INVX1 U29 ( .A(\write<7> ), .Y(n27) );
  INVX1 U30 ( .A(\write<8> ), .Y(n25) );
  INVX1 U31 ( .A(\write<9> ), .Y(n23) );
  INVX1 U32 ( .A(\write<10> ), .Y(n21) );
  INVX1 U33 ( .A(\write<12> ), .Y(n17) );
  INVX1 U34 ( .A(\write<13> ), .Y(n15) );
  INVX1 U35 ( .A(\write<14> ), .Y(n13) );
  INVX1 U36 ( .A(\write<15> ), .Y(n11) );
  INVX1 U37 ( .A(\write<11> ), .Y(n19) );
  INVX1 U38 ( .A(n3), .Y(n14) );
  INVX1 U39 ( .A(n4), .Y(n12) );
  BUFX2 U40 ( .A(\read<12> ), .Y(n5) );
  INVX1 U41 ( .A(n5), .Y(n18) );
  MUX2X1 U42 ( .B(n12), .A(n11), .S(n7), .Y(n57) );
  MUX2X1 U43 ( .B(n14), .A(n13), .S(n7), .Y(n56) );
  MUX2X1 U44 ( .B(n16), .A(n15), .S(n7), .Y(n55) );
  MUX2X1 U45 ( .B(n18), .A(n17), .S(n7), .Y(n54) );
  MUX2X1 U46 ( .B(n20), .A(n19), .S(n6), .Y(n53) );
  MUX2X1 U47 ( .B(n22), .A(n21), .S(n6), .Y(n52) );
  MUX2X1 U48 ( .B(n24), .A(n23), .S(n6), .Y(n51) );
  MUX2X1 U49 ( .B(n26), .A(n25), .S(n6), .Y(n50) );
  MUX2X1 U50 ( .B(n10), .A(n27), .S(n6), .Y(n49) );
  MUX2X1 U51 ( .B(n29), .A(n28), .S(n6), .Y(n48) );
  MUX2X1 U52 ( .B(n31), .A(n30), .S(n6), .Y(n47) );
  MUX2X1 U53 ( .B(n33), .A(n32), .S(n6), .Y(n46) );
  MUX2X1 U54 ( .B(n35), .A(n34), .S(n6), .Y(n45) );
  MUX2X1 U55 ( .B(n37), .A(n36), .S(n6), .Y(n44) );
  MUX2X1 U56 ( .B(n39), .A(n38), .S(n6), .Y(n43) );
  MUX2X1 U57 ( .B(n41), .A(n40), .S(n6), .Y(n42) );
endmodule


module reg16_32 ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51;

  dff_572 d0 ( .q(\read<0> ), .d(n36), .clk(clk), .rst(rst) );
  dff_571 d1 ( .q(\read<1> ), .d(n37), .clk(clk), .rst(rst) );
  dff_570 d2 ( .q(\read<2> ), .d(n38), .clk(clk), .rst(rst) );
  dff_569 d3 ( .q(\read<3> ), .d(n39), .clk(clk), .rst(rst) );
  dff_568 d4 ( .q(\read<4> ), .d(n40), .clk(clk), .rst(rst) );
  dff_567 d5 ( .q(\read<5> ), .d(n41), .clk(clk), .rst(rst) );
  dff_566 d6 ( .q(\read<6> ), .d(n42), .clk(clk), .rst(rst) );
  dff_565 d7 ( .q(\read<7> ), .d(n43), .clk(clk), .rst(rst) );
  dff_564 d8 ( .q(\read<8> ), .d(n44), .clk(clk), .rst(rst) );
  dff_563 d9 ( .q(\read<9> ), .d(n45), .clk(clk), .rst(rst) );
  dff_562 d10 ( .q(\read<10> ), .d(n46), .clk(clk), .rst(rst) );
  dff_561 d11 ( .q(\read<11> ), .d(n47), .clk(clk), .rst(rst) );
  dff_560 d12 ( .q(\read<12> ), .d(n48), .clk(clk), .rst(rst) );
  dff_559 d13 ( .q(\read<13> ), .d(n49), .clk(clk), .rst(rst) );
  dff_558 d14 ( .q(\read<14> ), .d(n50), .clk(clk), .rst(rst) );
  dff_557 d15 ( .q(\read<15> ), .d(n51), .clk(clk), .rst(rst) );
  INVX1 U1 ( .A(wr_en), .Y(n3) );
  INVX1 U2 ( .A(n3), .Y(n1) );
  INVX1 U3 ( .A(n3), .Y(n2) );
  INVX1 U4 ( .A(\read<0> ), .Y(n35) );
  INVX1 U5 ( .A(\read<1> ), .Y(n33) );
  INVX1 U6 ( .A(\read<2> ), .Y(n31) );
  INVX1 U7 ( .A(\read<3> ), .Y(n29) );
  INVX1 U8 ( .A(\read<4> ), .Y(n27) );
  INVX1 U9 ( .A(\read<5> ), .Y(n25) );
  INVX1 U10 ( .A(\read<6> ), .Y(n23) );
  INVX1 U11 ( .A(\read<7> ), .Y(n21) );
  INVX1 U12 ( .A(\read<8> ), .Y(n19) );
  INVX1 U13 ( .A(\read<9> ), .Y(n17) );
  INVX1 U14 ( .A(\read<10> ), .Y(n15) );
  INVX1 U15 ( .A(\read<11> ), .Y(n13) );
  INVX1 U16 ( .A(\read<12> ), .Y(n11) );
  INVX1 U17 ( .A(\read<13> ), .Y(n9) );
  INVX1 U18 ( .A(\read<14> ), .Y(n7) );
  INVX1 U19 ( .A(\read<15> ), .Y(n5) );
  INVX1 U20 ( .A(\write<0> ), .Y(n34) );
  INVX1 U21 ( .A(\write<1> ), .Y(n32) );
  INVX1 U22 ( .A(\write<2> ), .Y(n30) );
  INVX1 U23 ( .A(\write<3> ), .Y(n28) );
  INVX1 U24 ( .A(\write<4> ), .Y(n26) );
  INVX1 U25 ( .A(\write<5> ), .Y(n24) );
  INVX1 U26 ( .A(\write<6> ), .Y(n22) );
  INVX1 U27 ( .A(\write<7> ), .Y(n20) );
  INVX1 U28 ( .A(\write<8> ), .Y(n18) );
  INVX1 U29 ( .A(\write<9> ), .Y(n16) );
  INVX1 U30 ( .A(\write<10> ), .Y(n14) );
  INVX1 U31 ( .A(\write<11> ), .Y(n12) );
  INVX1 U32 ( .A(\write<12> ), .Y(n10) );
  INVX1 U33 ( .A(\write<13> ), .Y(n8) );
  INVX1 U34 ( .A(\write<14> ), .Y(n6) );
  INVX1 U35 ( .A(\write<15> ), .Y(n4) );
  MUX2X1 U36 ( .B(n5), .A(n4), .S(n2), .Y(n51) );
  MUX2X1 U37 ( .B(n7), .A(n6), .S(n2), .Y(n50) );
  MUX2X1 U38 ( .B(n9), .A(n8), .S(n2), .Y(n49) );
  MUX2X1 U39 ( .B(n11), .A(n10), .S(n2), .Y(n48) );
  MUX2X1 U40 ( .B(n13), .A(n12), .S(n1), .Y(n47) );
  MUX2X1 U41 ( .B(n15), .A(n14), .S(n1), .Y(n46) );
  MUX2X1 U42 ( .B(n17), .A(n16), .S(n1), .Y(n45) );
  MUX2X1 U43 ( .B(n19), .A(n18), .S(n1), .Y(n44) );
  MUX2X1 U44 ( .B(n21), .A(n20), .S(n1), .Y(n43) );
  MUX2X1 U45 ( .B(n23), .A(n22), .S(n1), .Y(n42) );
  MUX2X1 U46 ( .B(n25), .A(n24), .S(n1), .Y(n41) );
  MUX2X1 U47 ( .B(n27), .A(n26), .S(n1), .Y(n40) );
  MUX2X1 U48 ( .B(n29), .A(n28), .S(n1), .Y(n39) );
  MUX2X1 U49 ( .B(n31), .A(n30), .S(n1), .Y(n38) );
  MUX2X1 U50 ( .B(n33), .A(n32), .S(n1), .Y(n37) );
  MUX2X1 U51 ( .B(n35), .A(n34), .S(n1), .Y(n36) );
endmodule


module reg16_31 ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51;

  dff_556 d0 ( .q(\read<0> ), .d(n36), .clk(clk), .rst(rst) );
  dff_555 d1 ( .q(\read<1> ), .d(n37), .clk(clk), .rst(rst) );
  dff_554 d2 ( .q(\read<2> ), .d(n38), .clk(clk), .rst(rst) );
  dff_553 d3 ( .q(\read<3> ), .d(n39), .clk(clk), .rst(rst) );
  dff_552 d4 ( .q(\read<4> ), .d(n40), .clk(clk), .rst(rst) );
  dff_551 d5 ( .q(\read<5> ), .d(n41), .clk(clk), .rst(rst) );
  dff_550 d6 ( .q(\read<6> ), .d(n42), .clk(clk), .rst(rst) );
  dff_549 d7 ( .q(\read<7> ), .d(n43), .clk(clk), .rst(rst) );
  dff_548 d8 ( .q(\read<8> ), .d(n44), .clk(clk), .rst(rst) );
  dff_547 d9 ( .q(\read<9> ), .d(n45), .clk(clk), .rst(rst) );
  dff_546 d10 ( .q(\read<10> ), .d(n46), .clk(clk), .rst(rst) );
  dff_545 d11 ( .q(\read<11> ), .d(n47), .clk(clk), .rst(rst) );
  dff_544 d12 ( .q(\read<12> ), .d(n48), .clk(clk), .rst(rst) );
  dff_543 d13 ( .q(\read<13> ), .d(n49), .clk(clk), .rst(rst) );
  dff_542 d14 ( .q(\read<14> ), .d(n50), .clk(clk), .rst(rst) );
  dff_541 d15 ( .q(\read<15> ), .d(n51), .clk(clk), .rst(rst) );
  INVX1 U1 ( .A(wr_en), .Y(n3) );
  INVX1 U2 ( .A(n3), .Y(n1) );
  INVX1 U3 ( .A(n3), .Y(n2) );
  INVX1 U4 ( .A(\read<0> ), .Y(n35) );
  INVX1 U5 ( .A(\read<1> ), .Y(n33) );
  INVX1 U6 ( .A(\read<2> ), .Y(n31) );
  INVX1 U7 ( .A(\read<3> ), .Y(n29) );
  INVX1 U8 ( .A(\read<4> ), .Y(n27) );
  INVX1 U9 ( .A(\read<5> ), .Y(n25) );
  INVX1 U10 ( .A(\read<6> ), .Y(n23) );
  INVX1 U11 ( .A(\read<7> ), .Y(n21) );
  INVX1 U12 ( .A(\read<8> ), .Y(n19) );
  INVX1 U13 ( .A(\read<9> ), .Y(n17) );
  INVX1 U14 ( .A(\read<10> ), .Y(n15) );
  INVX1 U15 ( .A(\read<11> ), .Y(n13) );
  INVX1 U16 ( .A(\read<12> ), .Y(n11) );
  INVX1 U17 ( .A(\read<13> ), .Y(n9) );
  INVX1 U18 ( .A(\read<14> ), .Y(n7) );
  INVX1 U19 ( .A(\read<15> ), .Y(n5) );
  INVX1 U20 ( .A(\write<0> ), .Y(n34) );
  INVX1 U21 ( .A(\write<1> ), .Y(n32) );
  INVX1 U22 ( .A(\write<2> ), .Y(n30) );
  INVX1 U23 ( .A(\write<3> ), .Y(n28) );
  INVX1 U24 ( .A(\write<4> ), .Y(n26) );
  INVX1 U25 ( .A(\write<5> ), .Y(n24) );
  INVX1 U26 ( .A(\write<6> ), .Y(n22) );
  INVX1 U27 ( .A(\write<7> ), .Y(n20) );
  INVX1 U28 ( .A(\write<8> ), .Y(n18) );
  INVX1 U29 ( .A(\write<9> ), .Y(n16) );
  INVX1 U30 ( .A(\write<10> ), .Y(n14) );
  INVX1 U31 ( .A(\write<11> ), .Y(n12) );
  INVX1 U32 ( .A(\write<12> ), .Y(n10) );
  INVX1 U33 ( .A(\write<13> ), .Y(n8) );
  INVX1 U34 ( .A(\write<14> ), .Y(n6) );
  INVX1 U35 ( .A(\write<15> ), .Y(n4) );
  MUX2X1 U36 ( .B(n5), .A(n4), .S(n2), .Y(n51) );
  MUX2X1 U37 ( .B(n7), .A(n6), .S(n2), .Y(n50) );
  MUX2X1 U38 ( .B(n9), .A(n8), .S(n2), .Y(n49) );
  MUX2X1 U39 ( .B(n11), .A(n10), .S(n2), .Y(n48) );
  MUX2X1 U40 ( .B(n13), .A(n12), .S(n1), .Y(n47) );
  MUX2X1 U41 ( .B(n15), .A(n14), .S(n1), .Y(n46) );
  MUX2X1 U42 ( .B(n17), .A(n16), .S(n1), .Y(n45) );
  MUX2X1 U43 ( .B(n19), .A(n18), .S(n1), .Y(n44) );
  MUX2X1 U44 ( .B(n21), .A(n20), .S(n1), .Y(n43) );
  MUX2X1 U45 ( .B(n23), .A(n22), .S(n1), .Y(n42) );
  MUX2X1 U46 ( .B(n25), .A(n24), .S(n1), .Y(n41) );
  MUX2X1 U47 ( .B(n27), .A(n26), .S(n1), .Y(n40) );
  MUX2X1 U48 ( .B(n29), .A(n28), .S(n1), .Y(n39) );
  MUX2X1 U49 ( .B(n31), .A(n30), .S(n1), .Y(n38) );
  MUX2X1 U50 ( .B(n33), .A(n32), .S(n1), .Y(n37) );
  MUX2X1 U51 ( .B(n35), .A(n34), .S(n1), .Y(n36) );
endmodule


module reg16_30 ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51;

  dff_540 d0 ( .q(\read<0> ), .d(n36), .clk(clk), .rst(rst) );
  dff_539 d1 ( .q(\read<1> ), .d(n37), .clk(clk), .rst(rst) );
  dff_538 d2 ( .q(\read<2> ), .d(n38), .clk(clk), .rst(rst) );
  dff_537 d3 ( .q(\read<3> ), .d(n39), .clk(clk), .rst(rst) );
  dff_536 d4 ( .q(\read<4> ), .d(n40), .clk(clk), .rst(rst) );
  dff_535 d5 ( .q(\read<5> ), .d(n41), .clk(clk), .rst(rst) );
  dff_534 d6 ( .q(\read<6> ), .d(n42), .clk(clk), .rst(rst) );
  dff_533 d7 ( .q(\read<7> ), .d(n43), .clk(clk), .rst(rst) );
  dff_532 d8 ( .q(\read<8> ), .d(n44), .clk(clk), .rst(rst) );
  dff_531 d9 ( .q(\read<9> ), .d(n45), .clk(clk), .rst(rst) );
  dff_530 d10 ( .q(\read<10> ), .d(n46), .clk(clk), .rst(rst) );
  dff_529 d11 ( .q(\read<11> ), .d(n47), .clk(clk), .rst(rst) );
  dff_528 d12 ( .q(\read<12> ), .d(n48), .clk(clk), .rst(rst) );
  dff_527 d13 ( .q(\read<13> ), .d(n49), .clk(clk), .rst(rst) );
  dff_526 d14 ( .q(\read<14> ), .d(n50), .clk(clk), .rst(rst) );
  dff_525 d15 ( .q(\read<15> ), .d(n51), .clk(clk), .rst(rst) );
  INVX1 U1 ( .A(wr_en), .Y(n3) );
  INVX1 U2 ( .A(n3), .Y(n1) );
  INVX1 U3 ( .A(n3), .Y(n2) );
  INVX1 U4 ( .A(\read<0> ), .Y(n35) );
  INVX1 U5 ( .A(\read<1> ), .Y(n33) );
  INVX1 U6 ( .A(\read<2> ), .Y(n31) );
  INVX1 U7 ( .A(\read<3> ), .Y(n29) );
  INVX1 U8 ( .A(\read<4> ), .Y(n27) );
  INVX1 U9 ( .A(\read<5> ), .Y(n25) );
  INVX1 U10 ( .A(\read<6> ), .Y(n23) );
  INVX1 U11 ( .A(\read<7> ), .Y(n21) );
  INVX1 U12 ( .A(\read<8> ), .Y(n19) );
  INVX1 U13 ( .A(\read<9> ), .Y(n17) );
  INVX1 U14 ( .A(\read<10> ), .Y(n15) );
  INVX1 U15 ( .A(\read<11> ), .Y(n13) );
  INVX1 U16 ( .A(\read<12> ), .Y(n11) );
  INVX1 U17 ( .A(\read<13> ), .Y(n9) );
  INVX1 U18 ( .A(\read<14> ), .Y(n7) );
  INVX1 U19 ( .A(\read<15> ), .Y(n5) );
  INVX1 U20 ( .A(\write<0> ), .Y(n34) );
  INVX1 U21 ( .A(\write<1> ), .Y(n32) );
  INVX1 U22 ( .A(\write<2> ), .Y(n30) );
  INVX1 U23 ( .A(\write<3> ), .Y(n28) );
  INVX1 U24 ( .A(\write<4> ), .Y(n26) );
  INVX1 U25 ( .A(\write<5> ), .Y(n24) );
  INVX1 U26 ( .A(\write<6> ), .Y(n22) );
  INVX1 U27 ( .A(\write<7> ), .Y(n20) );
  INVX1 U28 ( .A(\write<8> ), .Y(n18) );
  INVX1 U29 ( .A(\write<9> ), .Y(n16) );
  INVX1 U30 ( .A(\write<10> ), .Y(n14) );
  INVX1 U31 ( .A(\write<11> ), .Y(n12) );
  INVX1 U32 ( .A(\write<12> ), .Y(n10) );
  INVX1 U33 ( .A(\write<13> ), .Y(n8) );
  INVX1 U34 ( .A(\write<14> ), .Y(n6) );
  INVX1 U35 ( .A(\write<15> ), .Y(n4) );
  MUX2X1 U36 ( .B(n5), .A(n4), .S(n2), .Y(n51) );
  MUX2X1 U37 ( .B(n7), .A(n6), .S(n2), .Y(n50) );
  MUX2X1 U38 ( .B(n9), .A(n8), .S(n2), .Y(n49) );
  MUX2X1 U39 ( .B(n11), .A(n10), .S(n2), .Y(n48) );
  MUX2X1 U40 ( .B(n13), .A(n12), .S(n1), .Y(n47) );
  MUX2X1 U41 ( .B(n15), .A(n14), .S(n1), .Y(n46) );
  MUX2X1 U42 ( .B(n17), .A(n16), .S(n1), .Y(n45) );
  MUX2X1 U43 ( .B(n19), .A(n18), .S(n1), .Y(n44) );
  MUX2X1 U44 ( .B(n21), .A(n20), .S(n1), .Y(n43) );
  MUX2X1 U45 ( .B(n23), .A(n22), .S(n1), .Y(n42) );
  MUX2X1 U46 ( .B(n25), .A(n24), .S(n1), .Y(n41) );
  MUX2X1 U47 ( .B(n27), .A(n26), .S(n1), .Y(n40) );
  MUX2X1 U48 ( .B(n29), .A(n28), .S(n1), .Y(n39) );
  MUX2X1 U49 ( .B(n31), .A(n30), .S(n1), .Y(n38) );
  MUX2X1 U50 ( .B(n33), .A(n32), .S(n1), .Y(n37) );
  MUX2X1 U51 ( .B(n35), .A(n34), .S(n1), .Y(n36) );
endmodule


module reg16_29 ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48;

  dff_524 d0 ( .q(\read<0> ), .d(n33), .clk(clk), .rst(rst) );
  dff_523 d1 ( .q(\read<1> ), .d(n34), .clk(clk), .rst(rst) );
  dff_522 d2 ( .q(\read<2> ), .d(n35), .clk(clk), .rst(rst) );
  dff_521 d3 ( .q(\read<3> ), .d(n36), .clk(clk), .rst(rst) );
  dff_520 d4 ( .q(\read<4> ), .d(n37), .clk(clk), .rst(rst) );
  dff_519 d5 ( .q(\read<5> ), .d(n38), .clk(clk), .rst(rst) );
  dff_518 d6 ( .q(\read<6> ), .d(n39), .clk(clk), .rst(rst) );
  dff_517 d7 ( .q(\read<7> ), .d(n40), .clk(clk), .rst(rst) );
  dff_516 d8 ( .q(\read<8> ), .d(n41), .clk(clk), .rst(rst) );
  dff_515 d9 ( .q(\read<9> ), .d(n42), .clk(clk), .rst(rst) );
  dff_514 d10 ( .q(\read<10> ), .d(n43), .clk(clk), .rst(rst) );
  dff_513 d11 ( .q(\read<11> ), .d(n44), .clk(clk), .rst(rst) );
  dff_512 d12 ( .q(\read<12> ), .d(n45), .clk(clk), .rst(rst) );
  dff_511 d13 ( .q(\read<13> ), .d(n46), .clk(clk), .rst(rst) );
  dff_510 d14 ( .q(\read<14> ), .d(n47), .clk(clk), .rst(rst) );
  dff_509 d15 ( .q(\read<15> ), .d(n48), .clk(clk), .rst(rst) );
  INVX1 U1 ( .A(\read<11> ), .Y(n10) );
  INVX1 U2 ( .A(\read<12> ), .Y(n8) );
  INVX1 U3 ( .A(\read<13> ), .Y(n6) );
  INVX1 U4 ( .A(\read<14> ), .Y(n4) );
  INVX1 U5 ( .A(\read<15> ), .Y(n2) );
  INVX1 U6 ( .A(\read<0> ), .Y(n32) );
  INVX1 U7 ( .A(\read<1> ), .Y(n30) );
  INVX1 U8 ( .A(\read<2> ), .Y(n28) );
  INVX1 U9 ( .A(\read<3> ), .Y(n26) );
  INVX1 U10 ( .A(\read<4> ), .Y(n24) );
  INVX1 U11 ( .A(\read<5> ), .Y(n22) );
  INVX1 U12 ( .A(\read<6> ), .Y(n20) );
  INVX1 U13 ( .A(\read<7> ), .Y(n18) );
  INVX1 U14 ( .A(\read<8> ), .Y(n16) );
  INVX1 U15 ( .A(\read<9> ), .Y(n14) );
  INVX1 U16 ( .A(\read<10> ), .Y(n12) );
  INVX1 U17 ( .A(\write<11> ), .Y(n9) );
  INVX1 U18 ( .A(\write<12> ), .Y(n7) );
  INVX1 U19 ( .A(\write<13> ), .Y(n5) );
  INVX1 U20 ( .A(\write<14> ), .Y(n3) );
  INVX1 U21 ( .A(\write<15> ), .Y(n1) );
  INVX1 U22 ( .A(\write<0> ), .Y(n31) );
  INVX1 U23 ( .A(\write<1> ), .Y(n29) );
  INVX1 U24 ( .A(\write<2> ), .Y(n27) );
  INVX1 U25 ( .A(\write<3> ), .Y(n25) );
  INVX1 U26 ( .A(\write<4> ), .Y(n23) );
  INVX1 U27 ( .A(\write<5> ), .Y(n21) );
  INVX1 U28 ( .A(\write<6> ), .Y(n19) );
  INVX1 U29 ( .A(\write<7> ), .Y(n17) );
  INVX1 U30 ( .A(\write<8> ), .Y(n15) );
  INVX1 U31 ( .A(\write<9> ), .Y(n13) );
  INVX1 U32 ( .A(\write<10> ), .Y(n11) );
  MUX2X1 U33 ( .B(n2), .A(n1), .S(wr_en), .Y(n48) );
  MUX2X1 U34 ( .B(n4), .A(n3), .S(wr_en), .Y(n47) );
  MUX2X1 U35 ( .B(n6), .A(n5), .S(wr_en), .Y(n46) );
  MUX2X1 U36 ( .B(n8), .A(n7), .S(wr_en), .Y(n45) );
  MUX2X1 U37 ( .B(n10), .A(n9), .S(wr_en), .Y(n44) );
  MUX2X1 U38 ( .B(n12), .A(n11), .S(wr_en), .Y(n43) );
  MUX2X1 U39 ( .B(n14), .A(n13), .S(wr_en), .Y(n42) );
  MUX2X1 U40 ( .B(n16), .A(n15), .S(wr_en), .Y(n41) );
  MUX2X1 U41 ( .B(n18), .A(n17), .S(wr_en), .Y(n40) );
  MUX2X1 U42 ( .B(n20), .A(n19), .S(wr_en), .Y(n39) );
  MUX2X1 U43 ( .B(n22), .A(n21), .S(wr_en), .Y(n38) );
  MUX2X1 U44 ( .B(n24), .A(n23), .S(wr_en), .Y(n37) );
  MUX2X1 U45 ( .B(n26), .A(n25), .S(wr_en), .Y(n36) );
  MUX2X1 U46 ( .B(n28), .A(n27), .S(wr_en), .Y(n35) );
  MUX2X1 U47 ( .B(n30), .A(n29), .S(wr_en), .Y(n34) );
  MUX2X1 U48 ( .B(n32), .A(n31), .S(wr_en), .Y(n33) );
endmodule


module reg1_23 ( d, q, clk, rst, en );
  input d, clk, rst, en;
  output q;
  wire   n1, n2, n3;

  dff_508 d0 ( .q(q), .d(n3), .clk(clk), .rst(rst) );
  INVX1 U1 ( .A(q), .Y(n2) );
  INVX1 U2 ( .A(d), .Y(n1) );
  MUX2X1 U3 ( .B(n2), .A(n1), .S(en), .Y(n3) );
endmodule


module reg1_22 ( d, q, clk, rst, en );
  input d, clk, rst, en;
  output q;
  wire   n1, n2, n3;

  dff_507 d0 ( .q(q), .d(n3), .clk(clk), .rst(rst) );
  INVX1 U1 ( .A(q), .Y(n2) );
  INVX1 U2 ( .A(d), .Y(n1) );
  MUX2X1 U3 ( .B(n2), .A(n1), .S(en), .Y(n3) );
endmodule


module reg16_28 ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48;

  dff_506 d0 ( .q(\read<0> ), .d(n33), .clk(clk), .rst(rst) );
  dff_505 d1 ( .q(\read<1> ), .d(n34), .clk(clk), .rst(rst) );
  dff_504 d2 ( .q(\read<2> ), .d(n35), .clk(clk), .rst(rst) );
  dff_503 d3 ( .q(\read<3> ), .d(n36), .clk(clk), .rst(rst) );
  dff_502 d4 ( .q(\read<4> ), .d(n37), .clk(clk), .rst(rst) );
  dff_501 d5 ( .q(\read<5> ), .d(n38), .clk(clk), .rst(rst) );
  dff_500 d6 ( .q(\read<6> ), .d(n39), .clk(clk), .rst(rst) );
  dff_499 d7 ( .q(\read<7> ), .d(n40), .clk(clk), .rst(rst) );
  dff_498 d8 ( .q(\read<8> ), .d(n41), .clk(clk), .rst(rst) );
  dff_497 d9 ( .q(\read<9> ), .d(n42), .clk(clk), .rst(rst) );
  dff_496 d10 ( .q(\read<10> ), .d(n43), .clk(clk), .rst(rst) );
  dff_495 d11 ( .q(\read<11> ), .d(n44), .clk(clk), .rst(rst) );
  dff_494 d12 ( .q(\read<12> ), .d(n45), .clk(clk), .rst(rst) );
  dff_493 d13 ( .q(\read<13> ), .d(n46), .clk(clk), .rst(rst) );
  dff_492 d14 ( .q(\read<14> ), .d(n47), .clk(clk), .rst(rst) );
  dff_491 d15 ( .q(\read<15> ), .d(n48), .clk(clk), .rst(rst) );
  INVX1 U1 ( .A(\read<0> ), .Y(n32) );
  INVX1 U2 ( .A(\read<1> ), .Y(n30) );
  INVX1 U3 ( .A(\read<2> ), .Y(n28) );
  INVX1 U4 ( .A(\read<3> ), .Y(n26) );
  INVX1 U5 ( .A(\read<4> ), .Y(n24) );
  INVX1 U6 ( .A(\read<5> ), .Y(n22) );
  INVX1 U7 ( .A(\read<6> ), .Y(n20) );
  INVX1 U8 ( .A(\read<7> ), .Y(n18) );
  INVX1 U9 ( .A(\read<8> ), .Y(n16) );
  INVX1 U10 ( .A(\read<9> ), .Y(n14) );
  INVX1 U11 ( .A(\read<10> ), .Y(n12) );
  INVX1 U12 ( .A(\read<11> ), .Y(n10) );
  INVX1 U13 ( .A(\read<12> ), .Y(n8) );
  INVX1 U14 ( .A(\read<13> ), .Y(n6) );
  INVX1 U15 ( .A(\read<14> ), .Y(n4) );
  INVX1 U16 ( .A(\read<15> ), .Y(n2) );
  INVX1 U17 ( .A(\write<0> ), .Y(n31) );
  INVX1 U18 ( .A(\write<1> ), .Y(n29) );
  INVX1 U19 ( .A(\write<2> ), .Y(n27) );
  INVX1 U20 ( .A(\write<3> ), .Y(n25) );
  INVX1 U21 ( .A(\write<4> ), .Y(n23) );
  INVX1 U22 ( .A(\write<5> ), .Y(n21) );
  INVX1 U23 ( .A(\write<6> ), .Y(n19) );
  INVX1 U24 ( .A(\write<7> ), .Y(n17) );
  INVX1 U25 ( .A(\write<8> ), .Y(n15) );
  INVX1 U26 ( .A(\write<9> ), .Y(n13) );
  INVX1 U27 ( .A(\write<10> ), .Y(n11) );
  INVX1 U28 ( .A(\write<11> ), .Y(n9) );
  INVX1 U29 ( .A(\write<12> ), .Y(n7) );
  INVX1 U30 ( .A(\write<13> ), .Y(n5) );
  INVX1 U31 ( .A(\write<14> ), .Y(n3) );
  INVX1 U32 ( .A(\write<15> ), .Y(n1) );
  MUX2X1 U33 ( .B(n2), .A(n1), .S(wr_en), .Y(n48) );
  MUX2X1 U34 ( .B(n4), .A(n3), .S(wr_en), .Y(n47) );
  MUX2X1 U35 ( .B(n6), .A(n5), .S(wr_en), .Y(n46) );
  MUX2X1 U36 ( .B(n8), .A(n7), .S(wr_en), .Y(n45) );
  MUX2X1 U37 ( .B(n10), .A(n9), .S(wr_en), .Y(n44) );
  MUX2X1 U38 ( .B(n12), .A(n11), .S(wr_en), .Y(n43) );
  MUX2X1 U39 ( .B(n14), .A(n13), .S(wr_en), .Y(n42) );
  MUX2X1 U40 ( .B(n16), .A(n15), .S(wr_en), .Y(n41) );
  MUX2X1 U41 ( .B(n18), .A(n17), .S(wr_en), .Y(n40) );
  MUX2X1 U42 ( .B(n20), .A(n19), .S(wr_en), .Y(n39) );
  MUX2X1 U43 ( .B(n22), .A(n21), .S(wr_en), .Y(n38) );
  MUX2X1 U44 ( .B(n24), .A(n23), .S(wr_en), .Y(n37) );
  MUX2X1 U45 ( .B(n26), .A(n25), .S(wr_en), .Y(n36) );
  MUX2X1 U46 ( .B(n28), .A(n27), .S(wr_en), .Y(n35) );
  MUX2X1 U47 ( .B(n30), .A(n29), .S(wr_en), .Y(n34) );
  MUX2X1 U48 ( .B(n32), .A(n31), .S(wr_en), .Y(n33) );
endmodule


module reg1_21 ( d, q, clk, rst, en );
  input d, clk, rst, en;
  output q;
  wire   n1, n2, n3;

  dff_490 d0 ( .q(q), .d(n3), .clk(clk), .rst(rst) );
  INVX1 U1 ( .A(q), .Y(n2) );
  INVX1 U2 ( .A(d), .Y(n1) );
  MUX2X1 U3 ( .B(n2), .A(n1), .S(en), .Y(n3) );
endmodule


module reg1_20 ( d, q, clk, rst, en );
  input d, clk, rst, en;
  output q;
  wire   n1, n2, n3;

  dff_489 d0 ( .q(q), .d(n3), .clk(clk), .rst(rst) );
  INVX1 U1 ( .A(q), .Y(n2) );
  INVX1 U2 ( .A(d), .Y(n1) );
  MUX2X1 U3 ( .B(n2), .A(n1), .S(en), .Y(n3) );
endmodule


module reg1_19 ( d, q, clk, rst, en );
  input d, clk, rst, en;
  output q;
  wire   n1, n2, n3;

  dff_488 d0 ( .q(q), .d(n3), .clk(clk), .rst(rst) );
  INVX1 U1 ( .A(q), .Y(n2) );
  INVX1 U2 ( .A(d), .Y(n1) );
  MUX2X1 U3 ( .B(n2), .A(n1), .S(en), .Y(n3) );
endmodule


module reg1_18 ( d, q, clk, rst, en );
  input d, clk, rst, en;
  output q;
  wire   n1, n2, n3;

  dff_487 d0 ( .q(q), .d(n3), .clk(clk), .rst(rst) );
  INVX1 U1 ( .A(q), .Y(n2) );
  INVX1 U2 ( .A(d), .Y(n1) );
  MUX2X1 U3 ( .B(n2), .A(n1), .S(en), .Y(n3) );
endmodule


module reg1_17 ( d, q, clk, rst, en );
  input d, clk, rst, en;
  output q;
  wire   n1, n2, n3;

  dff_486 d0 ( .q(q), .d(n3), .clk(clk), .rst(rst) );
  INVX1 U1 ( .A(q), .Y(n2) );
  INVX1 U2 ( .A(d), .Y(n1) );
  MUX2X1 U3 ( .B(n2), .A(n1), .S(en), .Y(n3) );
endmodule


module reg16_27 ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48;

  dff_485 d0 ( .q(\read<0> ), .d(n33), .clk(clk), .rst(rst) );
  dff_484 d1 ( .q(\read<1> ), .d(n34), .clk(clk), .rst(rst) );
  dff_483 d2 ( .q(\read<2> ), .d(n35), .clk(clk), .rst(rst) );
  dff_482 d3 ( .q(\read<3> ), .d(n36), .clk(clk), .rst(rst) );
  dff_481 d4 ( .q(\read<4> ), .d(n37), .clk(clk), .rst(rst) );
  dff_480 d5 ( .q(\read<5> ), .d(n38), .clk(clk), .rst(rst) );
  dff_479 d6 ( .q(\read<6> ), .d(n39), .clk(clk), .rst(rst) );
  dff_478 d7 ( .q(\read<7> ), .d(n40), .clk(clk), .rst(rst) );
  dff_477 d8 ( .q(\read<8> ), .d(n41), .clk(clk), .rst(rst) );
  dff_476 d9 ( .q(\read<9> ), .d(n42), .clk(clk), .rst(rst) );
  dff_475 d10 ( .q(\read<10> ), .d(n43), .clk(clk), .rst(rst) );
  dff_474 d11 ( .q(\read<11> ), .d(n44), .clk(clk), .rst(rst) );
  dff_473 d12 ( .q(\read<12> ), .d(n45), .clk(clk), .rst(rst) );
  dff_472 d13 ( .q(\read<13> ), .d(n46), .clk(clk), .rst(rst) );
  dff_471 d14 ( .q(\read<14> ), .d(n47), .clk(clk), .rst(rst) );
  dff_470 d15 ( .q(\read<15> ), .d(n48), .clk(clk), .rst(rst) );
  INVX1 U1 ( .A(\read<0> ), .Y(n32) );
  INVX1 U2 ( .A(\read<1> ), .Y(n30) );
  INVX1 U3 ( .A(\read<2> ), .Y(n28) );
  INVX1 U4 ( .A(\read<3> ), .Y(n26) );
  INVX1 U5 ( .A(\read<4> ), .Y(n24) );
  INVX1 U6 ( .A(\read<5> ), .Y(n22) );
  INVX1 U7 ( .A(\read<6> ), .Y(n20) );
  INVX1 U8 ( .A(\read<7> ), .Y(n18) );
  INVX1 U9 ( .A(\read<8> ), .Y(n16) );
  INVX1 U10 ( .A(\read<9> ), .Y(n14) );
  INVX1 U11 ( .A(\read<10> ), .Y(n12) );
  INVX1 U12 ( .A(\read<11> ), .Y(n10) );
  INVX1 U13 ( .A(\read<12> ), .Y(n8) );
  INVX1 U14 ( .A(\read<13> ), .Y(n6) );
  INVX1 U15 ( .A(\read<14> ), .Y(n4) );
  INVX1 U16 ( .A(\read<15> ), .Y(n2) );
  INVX1 U17 ( .A(\write<0> ), .Y(n31) );
  INVX1 U18 ( .A(\write<1> ), .Y(n29) );
  INVX1 U19 ( .A(\write<2> ), .Y(n27) );
  INVX1 U20 ( .A(\write<3> ), .Y(n25) );
  INVX1 U21 ( .A(\write<4> ), .Y(n23) );
  INVX1 U22 ( .A(\write<5> ), .Y(n21) );
  INVX1 U23 ( .A(\write<6> ), .Y(n19) );
  INVX1 U24 ( .A(\write<7> ), .Y(n17) );
  INVX1 U25 ( .A(\write<8> ), .Y(n15) );
  INVX1 U26 ( .A(\write<9> ), .Y(n13) );
  INVX1 U27 ( .A(\write<10> ), .Y(n11) );
  INVX1 U28 ( .A(\write<11> ), .Y(n9) );
  INVX1 U29 ( .A(\write<12> ), .Y(n7) );
  INVX1 U30 ( .A(\write<13> ), .Y(n5) );
  INVX1 U31 ( .A(\write<14> ), .Y(n3) );
  INVX1 U32 ( .A(\write<15> ), .Y(n1) );
  MUX2X1 U33 ( .B(n2), .A(n1), .S(wr_en), .Y(n48) );
  MUX2X1 U34 ( .B(n4), .A(n3), .S(wr_en), .Y(n47) );
  MUX2X1 U35 ( .B(n6), .A(n5), .S(wr_en), .Y(n46) );
  MUX2X1 U36 ( .B(n8), .A(n7), .S(wr_en), .Y(n45) );
  MUX2X1 U37 ( .B(n10), .A(n9), .S(wr_en), .Y(n44) );
  MUX2X1 U38 ( .B(n12), .A(n11), .S(wr_en), .Y(n43) );
  MUX2X1 U39 ( .B(n14), .A(n13), .S(wr_en), .Y(n42) );
  MUX2X1 U40 ( .B(n16), .A(n15), .S(wr_en), .Y(n41) );
  MUX2X1 U41 ( .B(n18), .A(n17), .S(wr_en), .Y(n40) );
  MUX2X1 U42 ( .B(n20), .A(n19), .S(wr_en), .Y(n39) );
  MUX2X1 U43 ( .B(n22), .A(n21), .S(wr_en), .Y(n38) );
  MUX2X1 U44 ( .B(n24), .A(n23), .S(wr_en), .Y(n37) );
  MUX2X1 U45 ( .B(n26), .A(n25), .S(wr_en), .Y(n36) );
  MUX2X1 U46 ( .B(n28), .A(n27), .S(wr_en), .Y(n35) );
  MUX2X1 U47 ( .B(n30), .A(n29), .S(wr_en), .Y(n34) );
  MUX2X1 U48 ( .B(n32), .A(n31), .S(wr_en), .Y(n33) );
endmodule


module reg16_26 ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60;

  dff_469 d0 ( .q(\read<0> ), .d(n46), .clk(clk), .rst(rst) );
  dff_468 d1 ( .q(\read<1> ), .d(n47), .clk(clk), .rst(rst) );
  dff_467 d2 ( .q(\read<2> ), .d(n48), .clk(clk), .rst(rst) );
  dff_466 d3 ( .q(\read<3> ), .d(n49), .clk(clk), .rst(rst) );
  dff_465 d4 ( .q(\read<4> ), .d(n50), .clk(clk), .rst(rst) );
  dff_464 d5 ( .q(\read<5> ), .d(n51), .clk(clk), .rst(rst) );
  dff_463 d6 ( .q(\read<6> ), .d(n52), .clk(clk), .rst(rst) );
  dff_462 d7 ( .q(\read<7> ), .d(n53), .clk(clk), .rst(rst) );
  dff_461 d8 ( .q(\read<8> ), .d(n54), .clk(clk), .rst(rst) );
  dff_460 d9 ( .q(\read<9> ), .d(n55), .clk(clk), .rst(rst) );
  dff_459 d10 ( .q(\read<10> ), .d(n56), .clk(clk), .rst(rst) );
  dff_458 d11 ( .q(\read<11> ), .d(n1), .clk(clk), .rst(rst) );
  dff_457 d12 ( .q(\read<12> ), .d(n57), .clk(clk), .rst(rst) );
  dff_456 d13 ( .q(\read<13> ), .d(n58), .clk(clk), .rst(rst) );
  dff_455 d14 ( .q(\read<14> ), .d(n59), .clk(clk), .rst(rst) );
  dff_454 d15 ( .q(\read<15> ), .d(n60), .clk(clk), .rst(rst) );
  INVX1 U1 ( .A(n17), .Y(n5) );
  INVX1 U2 ( .A(n19), .Y(n17) );
  INVX1 U3 ( .A(n17), .Y(n7) );
  INVX1 U4 ( .A(n17), .Y(n4) );
  INVX1 U5 ( .A(\read<1> ), .Y(n43) );
  INVX1 U6 ( .A(n17), .Y(n6) );
  INVX1 U7 ( .A(\read<4> ), .Y(n37) );
  INVX1 U8 ( .A(n17), .Y(n13) );
  INVX1 U9 ( .A(\read<5> ), .Y(n35) );
  INVX1 U10 ( .A(n17), .Y(n14) );
  INVX1 U11 ( .A(\read<6> ), .Y(n33) );
  INVX1 U12 ( .A(n17), .Y(n12) );
  INVX1 U13 ( .A(\read<7> ), .Y(n31) );
  INVX1 U14 ( .A(n17), .Y(n11) );
  INVX1 U15 ( .A(\read<9> ), .Y(n29) );
  INVX1 U16 ( .A(\write<11> ), .Y(n3) );
  INVX1 U17 ( .A(wr_en), .Y(n19) );
  INVX1 U18 ( .A(\read<11> ), .Y(n2) );
  INVX1 U19 ( .A(\read<12> ), .Y(n27) );
  INVX1 U20 ( .A(n18), .Y(n15) );
  INVX1 U21 ( .A(\read<13> ), .Y(n25) );
  INVX1 U22 ( .A(n18), .Y(n16) );
  INVX1 U23 ( .A(\read<14> ), .Y(n23) );
  INVX1 U24 ( .A(\read<15> ), .Y(n21) );
  INVX1 U25 ( .A(\read<0> ), .Y(n45) );
  INVX1 U26 ( .A(\read<2> ), .Y(n41) );
  INVX1 U27 ( .A(\read<3> ), .Y(n39) );
  INVX1 U28 ( .A(n8), .Y(n54) );
  INVX1 U29 ( .A(n19), .Y(n18) );
  INVX1 U30 ( .A(n18), .Y(n10) );
  MUX2X1 U31 ( .B(n3), .A(n2), .S(n19), .Y(n1) );
  INVX1 U32 ( .A(n9), .Y(n56) );
  MUX2X1 U33 ( .B(n38), .A(n39), .S(n4), .Y(n49) );
  MUX2X1 U34 ( .B(n44), .A(n45), .S(n5), .Y(n46) );
  MUX2X1 U35 ( .B(n36), .A(n37), .S(n6), .Y(n50) );
  INVX1 U36 ( .A(\write<1> ), .Y(n42) );
  INVX1 U37 ( .A(\write<3> ), .Y(n38) );
  MUX2X1 U38 ( .B(n40), .A(n41), .S(n7), .Y(n48) );
  INVX1 U39 ( .A(\write<4> ), .Y(n36) );
  MUX2X1 U40 ( .B(\read<8> ), .A(\write<8> ), .S(n17), .Y(n8) );
  MUX2X1 U41 ( .B(\read<10> ), .A(\write<10> ), .S(n17), .Y(n9) );
  INVX1 U42 ( .A(\write<0> ), .Y(n44) );
  MUX2X1 U43 ( .B(n26), .A(n27), .S(n10), .Y(n57) );
  INVX1 U44 ( .A(\write<2> ), .Y(n40) );
  INVX1 U45 ( .A(\write<12> ), .Y(n26) );
  MUX2X1 U46 ( .B(n28), .A(n29), .S(n11), .Y(n55) );
  MUX2X1 U47 ( .B(n30), .A(n31), .S(n12), .Y(n53) );
  MUX2X1 U48 ( .B(n34), .A(n35), .S(n13), .Y(n51) );
  MUX2X1 U49 ( .B(n32), .A(n33), .S(n14), .Y(n52) );
  INVX1 U50 ( .A(\write<6> ), .Y(n32) );
  INVX1 U51 ( .A(\write<9> ), .Y(n28) );
  INVX1 U52 ( .A(\write<7> ), .Y(n30) );
  MUX2X1 U53 ( .B(n24), .A(n25), .S(n15), .Y(n58) );
  INVX1 U54 ( .A(\write<5> ), .Y(n34) );
  MUX2X1 U55 ( .B(n22), .A(n23), .S(n16), .Y(n59) );
  INVX1 U56 ( .A(\write<13> ), .Y(n24) );
  MUX2X1 U57 ( .B(n20), .A(n21), .S(n10), .Y(n60) );
  INVX1 U58 ( .A(\write<15> ), .Y(n20) );
  INVX1 U59 ( .A(\write<14> ), .Y(n22) );
  MUX2X1 U60 ( .B(n43), .A(n42), .S(n17), .Y(n47) );
endmodule


module reg1_16 ( d, q, clk, rst, en );
  input d, clk, rst, en;
  output q;
  wire   n1, n2, n3;

  dff_453 d0 ( .q(q), .d(n3), .clk(clk), .rst(rst) );
  INVX1 U1 ( .A(q), .Y(n2) );
  INVX1 U2 ( .A(d), .Y(n1) );
  MUX2X1 U3 ( .B(n2), .A(n1), .S(en), .Y(n3) );
endmodule


module reg1_15 ( d, q, clk, rst, en );
  input d, clk, rst, en;
  output q;
  wire   n1, n2, n3;

  dff_452 d0 ( .q(q), .d(n3), .clk(clk), .rst(rst) );
  INVX1 U1 ( .A(q), .Y(n2) );
  INVX1 U2 ( .A(d), .Y(n1) );
  MUX2X1 U3 ( .B(n2), .A(n1), .S(en), .Y(n3) );
endmodule


module EX_control ( .ALUOp({\ALUOp<4> , \ALUOp<3> , \ALUOp<2> , \ALUOp<1> , 
        \ALUOp<0> }), ALUSrc, wr_r7, compareS_EX, .opcode({\opcode<4> , 
        \opcode<3> , \opcode<2> , \opcode<1> , \opcode<0> }) );
  input \opcode<4> , \opcode<3> , \opcode<2> , \opcode<1> , \opcode<0> ;
  output \ALUOp<4> , \ALUOp<3> , \ALUOp<2> , \ALUOp<1> , \ALUOp<0> , ALUSrc,
         wr_r7, compareS_EX;
  wire   n5, n6, n9, n11, n1, n2, n3, n4, n7, n10, n12, n13, n14, n16, n18;
  assign compareS_EX = 1'b1;

  NAND2X1 U10 ( .A(n9), .B(n13), .Y(\ALUOp<1> ) );
  NAND3X1 U11 ( .A(\opcode<2> ), .B(\opcode<1> ), .C(n12), .Y(n6) );
  OAI21X1 U13 ( .A(\opcode<4> ), .B(\opcode<3> ), .C(\opcode<1> ), .Y(n9) );
  OAI21X1 U14 ( .A(n16), .B(n5), .C(n11), .Y(\ALUOp<0> ) );
  OAI21X1 U15 ( .A(\opcode<4> ), .B(\opcode<2> ), .C(\opcode<0> ), .Y(n11) );
  INVX1 U2 ( .A(n14), .Y(\ALUOp<2> ) );
  INVX1 U3 ( .A(n16), .Y(\ALUOp<3> ) );
  INVX1 U4 ( .A(n18), .Y(\ALUOp<4> ) );
  INVX1 U5 ( .A(n13), .Y(wr_r7) );
  INVX1 U6 ( .A(n7), .Y(ALUSrc) );
  INVX1 U7 ( .A(\opcode<2> ), .Y(n14) );
  INVX1 U8 ( .A(\opcode<0> ), .Y(n5) );
  OR2X2 U9 ( .A(\opcode<4> ), .B(\opcode<3> ), .Y(n10) );
  AND2X2 U12 ( .A(\opcode<4> ), .B(\opcode<3> ), .Y(n1) );
  INVX1 U16 ( .A(n1), .Y(n2) );
  OR2X2 U17 ( .A(\opcode<2> ), .B(\opcode<1> ), .Y(n3) );
  INVX1 U18 ( .A(n3), .Y(n4) );
  OR2X2 U19 ( .A(n4), .B(n2), .Y(n7) );
  INVX1 U20 ( .A(n10), .Y(n12) );
  BUFX2 U21 ( .A(n6), .Y(n13) );
  INVX1 U22 ( .A(\opcode<4> ), .Y(n18) );
  INVX1 U23 ( .A(\opcode<3> ), .Y(n16) );
endmodule


module alu ( .A({\A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> , 
        \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , \A<0> 
        }), .B({\B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , \B<9> , 
        \B<8> , \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , \B<0> 
        }), Cin, .Op({\Op<2> , \Op<1> , \Op<0> }), invA, invB, sign, .Out({
        \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> , 
        \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , 
        \Out<2> , \Out<1> , \Out<0> }), Ofl, Z, N, P, c_out );
  input \A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> , \A<8> ,
         \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , \A<0> ,
         \B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , \B<9> , \B<8> ,
         \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , \B<0> , Cin,
         \Op<2> , \Op<1> , \Op<0> , invA, invB, sign;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> , Ofl, Z, N, P, c_out;
  wire   \opB<15> , \shiftOut<15> , \shiftOut<14> , \shiftOut<13> ,
         \shiftOut<12> , \shiftOut<11> , \shiftOut<10> , \shiftOut<9> ,
         \shiftOut<8> , \shiftOut<7> , \shiftOut<6> , \shiftOut<5> ,
         \shiftOut<4> , \shiftOut<2> , \shiftOut<1> , \shiftOut<0> ,
         \sumOut<15> , \sumOut<14> , \sumOut<13> , \sumOut<12> , \sumOut<11> ,
         \sumOut<10> , \sumOut<9> , \sumOut<8> , \sumOut<7> , \sumOut<6> ,
         \sumOut<5> , \sumOut<4> , \sumOut<3> , \sumOut<2> , \sumOut<1> ,
         \sumOut<0> , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n114, n116, n118, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n262, n264, n266, n268, n270, n272, n274, n276,
         n278, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492;

  shifter shift ( .In({n324, n446, n467, n468, n323, n449, n457, n453, n452, 
        n450, n458, n448, n451, n318, n455, n454}), .Cnt({n456, n459, n460, 
        n73}), .Op({\Op<1> , \Op<0> }), .Out({\shiftOut<15> , \shiftOut<14> , 
        \shiftOut<13> , \shiftOut<12> , \shiftOut<11> , \shiftOut<10> , 
        \shiftOut<9> , \shiftOut<8> , \shiftOut<7> , \shiftOut<6> , 
        \shiftOut<5> , \shiftOut<4> , n461, \shiftOut<2> , \shiftOut<1> , 
        \shiftOut<0> }) );
  CLA16_0 adder ( .A({n13, n466, n467, n20, n469, n470, n471, n35, n472, n473, 
        n474, n475, n476, n477, n478, n479}), .B({\opB<15> , n480, n26, n481, 
        n482, n483, n65, n484, n485, n486, n487, n488, n489, n490, n491, n492}), .Cin(Cin), .Cout(c_out), .S({\sumOut<15> , \sumOut<14> , \sumOut<13> , 
        \sumOut<12> , \sumOut<11> , \sumOut<10> , \sumOut<9> , \sumOut<8> , 
        \sumOut<7> , \sumOut<6> , \sumOut<5> , \sumOut<4> , \sumOut<3> , 
        \sumOut<2> , \sumOut<1> , \sumOut<0> }) );
  BUFX2 U1 ( .A(n460), .Y(n1) );
  INVX1 U2 ( .A(n321), .Y(n490) );
  AND2X2 U3 ( .A(n195), .B(n132), .Y(n96) );
  INVX2 U4 ( .A(n362), .Y(n459) );
  INVX2 U5 ( .A(n347), .Y(n456) );
  INVX1 U6 ( .A(n1), .Y(n2) );
  OR2X2 U7 ( .A(n280), .B(n4), .Y(n3) );
  INVX8 U8 ( .A(n317), .Y(n4) );
  OR2X2 U9 ( .A(n198), .B(n6), .Y(n5) );
  INVX1 U10 ( .A(n5), .Y(n116) );
  INVX8 U11 ( .A(n438), .Y(n6) );
  INVX1 U12 ( .A(n362), .Y(n7) );
  XOR2X1 U13 ( .A(\B<2> ), .B(n8), .Y(n321) );
  INVX8 U14 ( .A(n42), .Y(n8) );
  OR2X2 U15 ( .A(n165), .B(n291), .Y(n9) );
  AND2X2 U16 ( .A(\sumOut<3> ), .B(n316), .Y(n291) );
  AND2X2 U17 ( .A(n79), .B(n100), .Y(n120) );
  INVX1 U18 ( .A(n74), .Y(n58) );
  INVX2 U19 ( .A(n14), .Y(n38) );
  INVX1 U20 ( .A(\opB<15> ), .Y(n49) );
  INVX1 U21 ( .A(n14), .Y(n29) );
  INVX1 U22 ( .A(n141), .Y(n343) );
  INVX2 U23 ( .A(n343), .Y(n342) );
  INVX2 U24 ( .A(n339), .Y(n21) );
  XOR2X1 U25 ( .A(n329), .B(n340), .Y(n10) );
  XOR2X1 U26 ( .A(n330), .B(n340), .Y(n11) );
  XOR2X1 U27 ( .A(\B<8> ), .B(n340), .Y(n12) );
  INVX2 U28 ( .A(n301), .Y(n344) );
  INVX1 U29 ( .A(n48), .Y(n435) );
  AND2X1 U30 ( .A(n316), .B(\sumOut<12> ), .Y(n285) );
  INVX1 U31 ( .A(n285), .Y(n37) );
  INVX2 U32 ( .A(n401), .Y(n457) );
  BUFX2 U33 ( .A(n324), .Y(n13) );
  INVX2 U34 ( .A(n70), .Y(n324) );
  XOR2X1 U35 ( .A(\B<14> ), .B(n42), .Y(n480) );
  XOR2X1 U36 ( .A(\A<4> ), .B(n14), .Y(n416) );
  INVX8 U37 ( .A(n341), .Y(n14) );
  BUFX2 U38 ( .A(n26), .Y(n15) );
  INVX4 U39 ( .A(n377), .Y(n454) );
  BUFX2 U40 ( .A(\shiftOut<11> ), .Y(n16) );
  BUFX2 U41 ( .A(n440), .Y(n17) );
  AND2X2 U42 ( .A(n312), .B(n313), .Y(n28) );
  INVX1 U43 ( .A(n145), .Y(n18) );
  INVX1 U44 ( .A(n454), .Y(n19) );
  BUFX2 U45 ( .A(n468), .Y(n20) );
  INVX2 U46 ( .A(n383), .Y(n468) );
  XNOR2X1 U47 ( .A(\A<10> ), .B(n14), .Y(n470) );
  XNOR2X1 U48 ( .A(\B<11> ), .B(n346), .Y(n482) );
  XOR2X1 U49 ( .A(\B<2> ), .B(n21), .Y(n362) );
  INVX1 U50 ( .A(\A<11> ), .Y(n22) );
  INVX1 U51 ( .A(n22), .Y(n23) );
  XOR2X1 U52 ( .A(n136), .B(n346), .Y(n492) );
  INVX1 U53 ( .A(n351), .Y(n453) );
  INVX1 U54 ( .A(n68), .Y(n24) );
  XNOR2X1 U55 ( .A(\A<0> ), .B(n14), .Y(n479) );
  AND2X2 U56 ( .A(\shiftOut<8> ), .B(n442), .Y(n304) );
  AND2X2 U57 ( .A(n118), .B(n440), .Y(n25) );
  INVX1 U58 ( .A(\sumOut<11> ), .Y(n72) );
  INVX2 U59 ( .A(n371), .Y(n446) );
  XOR2X1 U60 ( .A(n122), .B(n21), .Y(n428) );
  XNOR2X1 U61 ( .A(n121), .B(n120), .Y(P) );
  XNOR2X1 U62 ( .A(\B<9> ), .B(n21), .Y(n65) );
  AND2X2 U63 ( .A(\sumOut<11> ), .B(n316), .Y(n167) );
  XNOR2X1 U64 ( .A(n27), .B(n339), .Y(n26) );
  INVX1 U65 ( .A(n15), .Y(n410) );
  INVX1 U66 ( .A(\B<13> ), .Y(n27) );
  XOR2X1 U67 ( .A(\A<7> ), .B(n29), .Y(n472) );
  AND2X2 U68 ( .A(\sumOut<7> ), .B(n316), .Y(n82) );
  INVX1 U69 ( .A(n320), .Y(n30) );
  AND2X2 U70 ( .A(n30), .B(n44), .Y(n31) );
  AND2X2 U71 ( .A(n187), .B(n450), .Y(n172) );
  INVX1 U72 ( .A(n448), .Y(n32) );
  XOR2X1 U73 ( .A(n33), .B(n341), .Y(n389) );
  INVX1 U74 ( .A(\A<10> ), .Y(n33) );
  AND2X2 U75 ( .A(n389), .B(n342), .Y(n229) );
  INVX1 U76 ( .A(n284), .Y(n34) );
  INVX1 U77 ( .A(n351), .Y(n35) );
  AND2X2 U78 ( .A(n36), .B(n25), .Y(n52) );
  AND2X2 U79 ( .A(n298), .B(n37), .Y(n36) );
  INVX2 U80 ( .A(n428), .Y(n460) );
  INVX1 U81 ( .A(n71), .Y(n332) );
  XNOR2X1 U82 ( .A(n23), .B(n341), .Y(n56) );
  XOR2X1 U83 ( .A(\B<7> ), .B(n42), .Y(n485) );
  XOR2X1 U84 ( .A(\A<2> ), .B(n38), .Y(n477) );
  BUFX2 U85 ( .A(n448), .Y(n39) );
  BUFX2 U86 ( .A(n308), .Y(n40) );
  XOR2X1 U87 ( .A(n41), .B(n341), .Y(n377) );
  INVX1 U88 ( .A(\A<0> ), .Y(n41) );
  AND2X2 U89 ( .A(n19), .B(n141), .Y(n221) );
  AND2X2 U90 ( .A(n452), .B(n189), .Y(n176) );
  XOR2X1 U91 ( .A(\B<3> ), .B(n42), .Y(n489) );
  INVX8 U92 ( .A(n346), .Y(n42) );
  INVX1 U93 ( .A(n393), .Y(n54) );
  INVX4 U94 ( .A(n349), .Y(n450) );
  INVX1 U95 ( .A(n96), .Y(n45) );
  XOR2X1 U96 ( .A(n43), .B(n339), .Y(n345) );
  INVX1 U97 ( .A(\B<6> ), .Y(n43) );
  OAI21X1 U98 ( .A(n442), .B(n45), .C(n150), .Y(n44) );
  INVX1 U99 ( .A(n311), .Y(n46) );
  INVX1 U100 ( .A(n311), .Y(\Out<15> ) );
  AND2X2 U101 ( .A(\sumOut<13> ), .B(n316), .Y(n169) );
  XOR2X1 U102 ( .A(\A<3> ), .B(n47), .Y(n476) );
  INVX8 U103 ( .A(n14), .Y(n47) );
  AND2X2 U104 ( .A(\sumOut<1> ), .B(n316), .Y(n194) );
  NOR3X1 U105 ( .A(n70), .B(n49), .C(\sumOut<15> ), .Y(n48) );
  AND2X2 U106 ( .A(n31), .B(n149), .Y(n143) );
  AND2X2 U107 ( .A(n344), .B(n424), .Y(n193) );
  INVX1 U108 ( .A(n312), .Y(\Out<7> ) );
  AND2X2 U109 ( .A(\sumOut<15> ), .B(n316), .Y(n97) );
  AND2X2 U110 ( .A(n53), .B(n52), .Y(n51) );
  NOR3X1 U111 ( .A(n54), .B(n331), .C(n84), .Y(n53) );
  XNOR2X1 U112 ( .A(\B<3> ), .B(n340), .Y(n347) );
  AND2X2 U113 ( .A(n401), .B(n342), .Y(n235) );
  OR2X2 U114 ( .A(n125), .B(n153), .Y(n55) );
  INVX4 U115 ( .A(n389), .Y(n449) );
  INVX4 U116 ( .A(n56), .Y(n323) );
  AND2X2 U117 ( .A(n486), .B(n353), .Y(n157) );
  AND2X2 U118 ( .A(n383), .B(n342), .Y(n225) );
  AND2X2 U119 ( .A(n32), .B(n342), .Y(n245) );
  AND2X2 U120 ( .A(n409), .B(n342), .Y(n241) );
  INVX1 U121 ( .A(n136), .Y(n57) );
  XOR2X1 U122 ( .A(\B<0> ), .B(n58), .Y(n73) );
  INVX1 U123 ( .A(n60), .Y(n59) );
  INVX1 U124 ( .A(n2), .Y(n60) );
  INVX4 U125 ( .A(n409), .Y(n467) );
  INVX4 U126 ( .A(n416), .Y(n448) );
  AND2X2 U127 ( .A(n199), .B(n185), .Y(n147) );
  INVX1 U128 ( .A(n290), .Y(n61) );
  BUFX2 U129 ( .A(\shiftOut<1> ), .Y(n62) );
  INVX1 U130 ( .A(n435), .Y(n63) );
  XOR2X1 U131 ( .A(\B<9> ), .B(n339), .Y(n64) );
  AND2X2 U132 ( .A(n126), .B(n155), .Y(n289) );
  INVX1 U133 ( .A(n64), .Y(n402) );
  AND2X2 U134 ( .A(n435), .B(n283), .Y(n262) );
  AND2X2 U135 ( .A(n316), .B(\sumOut<9> ), .Y(n287) );
  AND2X2 U136 ( .A(\sumOut<10> ), .B(n316), .Y(n331) );
  INVX1 U137 ( .A(n313), .Y(\Out<6> ) );
  AND2X2 U138 ( .A(n323), .B(n191), .Y(n178) );
  AND2X2 U139 ( .A(n286), .B(n298), .Y(n272) );
  XNOR2X1 U140 ( .A(n57), .B(n74), .Y(n67) );
  INVX2 U141 ( .A(n339), .Y(n74) );
  NOR3X1 U142 ( .A(n290), .B(n296), .C(n18), .Y(n68) );
  INVX1 U143 ( .A(n122), .Y(n69) );
  XNOR2X1 U144 ( .A(n69), .B(n340), .Y(n491) );
  XNOR2X1 U145 ( .A(\A<15> ), .B(n341), .Y(n70) );
  AND2X2 U146 ( .A(n98), .B(n214), .Y(n311) );
  AND2X2 U147 ( .A(n297), .B(n61), .Y(n214) );
  AND2X2 U148 ( .A(\sumOut<5> ), .B(n316), .Y(n180) );
  AND2X2 U149 ( .A(n144), .B(n335), .Y(n264) );
  OAI21X1 U150 ( .A(n317), .B(n72), .C(n376), .Y(n71) );
  OR2X2 U151 ( .A(\shiftOut<11> ), .B(n315), .Y(n334) );
  AND2X2 U152 ( .A(\shiftOut<14> ), .B(n442), .Y(n125) );
  AND2X2 U153 ( .A(n37), .B(n289), .Y(n276) );
  OR2X2 U154 ( .A(n294), .B(n300), .Y(n75) );
  INVX1 U155 ( .A(n75), .Y(n76) );
  AND2X2 U156 ( .A(n111), .B(n143), .Y(n77) );
  AND2X2 U157 ( .A(n442), .B(\shiftOut<4> ), .Y(n165) );
  AND2X2 U158 ( .A(n336), .B(\Out<15> ), .Y(n78) );
  INVX1 U159 ( .A(n78), .Y(n79) );
  AND2X2 U160 ( .A(\sumOut<6> ), .B(n316), .Y(n80) );
  INVX1 U161 ( .A(n80), .Y(n81) );
  AND2X2 U162 ( .A(n442), .B(n109), .Y(n83) );
  OR2X2 U163 ( .A(n5), .B(n288), .Y(n84) );
  AND2X2 U164 ( .A(n134), .B(n442), .Y(n85) );
  INVX1 U165 ( .A(n85), .Y(n86) );
  AND2X2 U166 ( .A(n442), .B(n112), .Y(n87) );
  INVX1 U167 ( .A(n87), .Y(n88) );
  AND2X2 U168 ( .A(\shiftOut<13> ), .B(n442), .Y(n89) );
  INVX1 U169 ( .A(n89), .Y(n90) );
  AND2X2 U170 ( .A(n316), .B(\sumOut<4> ), .Y(n91) );
  AND2X2 U171 ( .A(n456), .B(n420), .Y(n92) );
  INVX1 U172 ( .A(n92), .Y(n93) );
  AND2X2 U173 ( .A(n344), .B(n426), .Y(n94) );
  INVX1 U174 ( .A(n94), .Y(n95) );
  INVX1 U175 ( .A(n97), .Y(n98) );
  AND2X2 U176 ( .A(n338), .B(n337), .Y(n99) );
  INVX1 U177 ( .A(n99), .Y(n100) );
  AND2X2 U178 ( .A(n442), .B(\shiftOut<2> ), .Y(n101) );
  INVX1 U179 ( .A(n101), .Y(n102) );
  AND2X2 U180 ( .A(n451), .B(n108), .Y(n103) );
  INVX1 U181 ( .A(n103), .Y(n104) );
  BUFX2 U182 ( .A(\shiftOut<0> ), .Y(n105) );
  BUFX2 U183 ( .A(n461), .Y(n106) );
  AND2X2 U184 ( .A(n344), .B(n421), .Y(n107) );
  INVX1 U185 ( .A(n107), .Y(n108) );
  BUFX2 U186 ( .A(\shiftOut<12> ), .Y(n109) );
  OR2X2 U187 ( .A(n9), .B(n304), .Y(n110) );
  INVX1 U188 ( .A(n110), .Y(n111) );
  BUFX2 U189 ( .A(\shiftOut<9> ), .Y(n112) );
  BUFX2 U190 ( .A(n462), .Y(\Out<3> ) );
  AND2X2 U191 ( .A(n96), .B(n140), .Y(n114) );
  INVX1 U192 ( .A(n114), .Y(\Out<1> ) );
  INVX1 U193 ( .A(n116), .Y(\Out<0> ) );
  AND2X2 U194 ( .A(n102), .B(n366), .Y(n118) );
  INVX1 U195 ( .A(n118), .Y(\Out<2> ) );
  BUFX2 U196 ( .A(n434), .Y(n121) );
  BUFX2 U197 ( .A(\B<1> ), .Y(n122) );
  INVX2 U198 ( .A(n348), .Y(n451) );
  INVX1 U199 ( .A(n180), .Y(n123) );
  INVX1 U200 ( .A(n82), .Y(n124) );
  INVX1 U201 ( .A(n83), .Y(n126) );
  INVX1 U202 ( .A(n356), .Y(n127) );
  INVX1 U203 ( .A(n127), .Y(n128) );
  AND2X2 U204 ( .A(n68), .B(n317), .Y(n129) );
  INVX1 U205 ( .A(n129), .Y(n130) );
  INVX1 U206 ( .A(n430), .Y(n131) );
  INVX1 U207 ( .A(n131), .Y(n132) );
  INVX1 U208 ( .A(\shiftOut<10> ), .Y(n133) );
  INVX1 U209 ( .A(n133), .Y(n134) );
  BUFX2 U210 ( .A(\B<5> ), .Y(n135) );
  INVX1 U211 ( .A(\B<0> ), .Y(n136) );
  AND2X2 U212 ( .A(n35), .B(n192), .Y(n137) );
  INVX1 U213 ( .A(n137), .Y(n138) );
  AND2X2 U214 ( .A(n62), .B(n442), .Y(n139) );
  INVX1 U215 ( .A(n139), .Y(n140) );
  INVX1 U216 ( .A(n422), .Y(n141) );
  INVX1 U217 ( .A(n141), .Y(n142) );
  AND2X1 U218 ( .A(\opB<15> ), .B(n406), .Y(n407) );
  AND2X2 U219 ( .A(n86), .B(n196), .Y(n144) );
  AND2X2 U220 ( .A(n90), .B(n197), .Y(n145) );
  INVX1 U221 ( .A(n145), .Y(n146) );
  OR2X2 U222 ( .A(n327), .B(n201), .Y(n148) );
  INVX1 U223 ( .A(n148), .Y(n149) );
  OR2X2 U224 ( .A(\shiftOut<1> ), .B(n295), .Y(n150) );
  INVX1 U225 ( .A(n359), .Y(n151) );
  INVX1 U226 ( .A(n151), .Y(n152) );
  INVX1 U227 ( .A(n154), .Y(n153) );
  BUFX2 U228 ( .A(n374), .Y(n154) );
  BUFX2 U229 ( .A(n386), .Y(n155) );
  BUFX2 U230 ( .A(n404), .Y(n156) );
  INVX1 U231 ( .A(n157), .Y(n158) );
  AND2X1 U232 ( .A(n10), .B(n357), .Y(n159) );
  INVX1 U233 ( .A(n159), .Y(n160) );
  AND2X1 U234 ( .A(n11), .B(n367), .Y(n161) );
  INVX1 U235 ( .A(n161), .Y(n162) );
  AND2X1 U236 ( .A(n12), .B(n423), .Y(n163) );
  INVX1 U237 ( .A(n163), .Y(n164) );
  INVX1 U238 ( .A(n165), .Y(n166) );
  INVX1 U239 ( .A(n167), .Y(n168) );
  INVX1 U240 ( .A(n169), .Y(n170) );
  BUFX2 U241 ( .A(n443), .Y(n171) );
  INVX1 U242 ( .A(n172), .Y(n173) );
  OR2X1 U243 ( .A(n442), .B(\Op<0> ), .Y(n174) );
  INVX1 U244 ( .A(n174), .Y(n175) );
  INVX1 U245 ( .A(n176), .Y(n177) );
  INVX1 U246 ( .A(n178), .Y(n179) );
  INVX1 U247 ( .A(n180), .Y(n181) );
  AND2X1 U248 ( .A(\sumOut<14> ), .B(n316), .Y(n182) );
  INVX1 U249 ( .A(n182), .Y(n183) );
  INVX1 U250 ( .A(n419), .Y(n184) );
  INVX1 U251 ( .A(n184), .Y(n185) );
  AND2X1 U252 ( .A(n344), .B(n354), .Y(n186) );
  INVX1 U253 ( .A(n186), .Y(n187) );
  AND2X1 U254 ( .A(n344), .B(n358), .Y(n188) );
  INVX1 U255 ( .A(n188), .Y(n189) );
  AND2X1 U256 ( .A(n344), .B(n368), .Y(n190) );
  INVX1 U257 ( .A(n190), .Y(n191) );
  INVX1 U258 ( .A(n193), .Y(n192) );
  INVX1 U259 ( .A(n194), .Y(n195) );
  BUFX2 U260 ( .A(n392), .Y(n196) );
  BUFX2 U261 ( .A(n412), .Y(n197) );
  AND2X2 U262 ( .A(n105), .B(n442), .Y(n198) );
  INVX1 U263 ( .A(n91), .Y(n199) );
  AND2X2 U264 ( .A(n147), .B(n76), .Y(n200) );
  INVX1 U265 ( .A(n200), .Y(n201) );
  BUFX2 U266 ( .A(n373), .Y(n202) );
  BUFX2 U267 ( .A(n385), .Y(n203) );
  BUFX2 U268 ( .A(n391), .Y(n204) );
  BUFX2 U269 ( .A(n403), .Y(n205) );
  BUFX2 U270 ( .A(n411), .Y(n206) );
  BUFX2 U271 ( .A(n418), .Y(n207) );
  INVX1 U272 ( .A(n429), .Y(n208) );
  INVX1 U273 ( .A(n208), .Y(n209) );
  AND2X2 U274 ( .A(n158), .B(n173), .Y(n210) );
  INVX1 U275 ( .A(n210), .Y(n211) );
  AND2X2 U276 ( .A(n160), .B(n177), .Y(n212) );
  INVX1 U277 ( .A(n212), .Y(n213) );
  INVX1 U278 ( .A(n146), .Y(n444) );
  AND2X1 U279 ( .A(n361), .B(n342), .Y(n215) );
  INVX1 U280 ( .A(n215), .Y(n216) );
  AND2X1 U281 ( .A(n344), .B(n370), .Y(n217) );
  INVX1 U282 ( .A(n217), .Y(n218) );
  AND2X2 U283 ( .A(n371), .B(n342), .Y(n219) );
  INVX1 U284 ( .A(n219), .Y(n220) );
  INVX1 U285 ( .A(n221), .Y(n222) );
  AND2X1 U286 ( .A(n344), .B(n382), .Y(n223) );
  INVX1 U287 ( .A(n223), .Y(n224) );
  INVX1 U288 ( .A(n225), .Y(n226) );
  AND2X1 U289 ( .A(n344), .B(n388), .Y(n227) );
  INVX1 U290 ( .A(n227), .Y(n228) );
  INVX1 U291 ( .A(n229), .Y(n230) );
  AND2X1 U292 ( .A(n395), .B(n342), .Y(n231) );
  INVX1 U293 ( .A(n231), .Y(n232) );
  AND2X1 U294 ( .A(n344), .B(n400), .Y(n233) );
  INVX1 U295 ( .A(n233), .Y(n234) );
  INVX1 U296 ( .A(n235), .Y(n236) );
  AND2X1 U297 ( .A(n344), .B(n405), .Y(n237) );
  INVX1 U298 ( .A(n237), .Y(n238) );
  AND2X1 U299 ( .A(n344), .B(n408), .Y(n239) );
  INVX1 U300 ( .A(n239), .Y(n240) );
  INVX1 U301 ( .A(n241), .Y(n242) );
  AND2X1 U302 ( .A(n344), .B(n415), .Y(n243) );
  INVX1 U303 ( .A(n243), .Y(n244) );
  INVX1 U304 ( .A(n245), .Y(n246) );
  AND2X1 U305 ( .A(n427), .B(n342), .Y(n247) );
  INVX1 U306 ( .A(n247), .Y(n248) );
  INVX1 U307 ( .A(n365), .Y(n249) );
  INVX1 U308 ( .A(n249), .Y(n250) );
  BUFX2 U309 ( .A(n397), .Y(n251) );
  INVX1 U310 ( .A(n364), .Y(n252) );
  INVX1 U311 ( .A(n252), .Y(n253) );
  INVX1 U312 ( .A(n380), .Y(n254) );
  INVX1 U313 ( .A(n254), .Y(n255) );
  BUFX2 U314 ( .A(n398), .Y(n256) );
  BUFX2 U315 ( .A(n379), .Y(n257) );
  INVX1 U316 ( .A(n77), .Y(n258) );
  AND2X1 U317 ( .A(\Op<0> ), .B(\Op<2> ), .Y(n259) );
  INVX1 U318 ( .A(n259), .Y(n260) );
  BUFX2 U319 ( .A(n447), .Y(\Out<8> ) );
  INVX1 U320 ( .A(n262), .Y(Ofl) );
  INVX1 U321 ( .A(n264), .Y(\Out<10> ) );
  AND2X2 U322 ( .A(n170), .B(n444), .Y(n266) );
  INVX1 U323 ( .A(n266), .Y(\Out<13> ) );
  AND2X2 U324 ( .A(n166), .B(n147), .Y(n268) );
  INVX1 U325 ( .A(n268), .Y(\Out<4> ) );
  AND2X2 U326 ( .A(n17), .B(n181), .Y(n270) );
  INVX1 U327 ( .A(n270), .Y(\Out<5> ) );
  INVX1 U328 ( .A(n272), .Y(\Out<9> ) );
  AND2X2 U329 ( .A(n168), .B(n171), .Y(n274) );
  INVX1 U330 ( .A(n274), .Y(\Out<11> ) );
  INVX1 U331 ( .A(n276), .Y(\Out<12> ) );
  AND2X2 U332 ( .A(n445), .B(n183), .Y(n278) );
  INVX1 U333 ( .A(n278), .Y(\Out<14> ) );
  INVX1 U334 ( .A(n333), .Y(n280) );
  INVX1 U335 ( .A(n280), .Y(n281) );
  INVX1 U336 ( .A(n284), .Y(n282) );
  INVX1 U337 ( .A(n282), .Y(n283) );
  BUFX2 U338 ( .A(n436), .Y(n284) );
  INVX1 U339 ( .A(n287), .Y(n286) );
  INVX1 U340 ( .A(n289), .Y(n288) );
  AND2X2 U341 ( .A(\shiftOut<15> ), .B(n442), .Y(n290) );
  INVX1 U342 ( .A(n291), .Y(n292) );
  AND2X2 U343 ( .A(n104), .B(n93), .Y(n293) );
  INVX1 U344 ( .A(n293), .Y(n294) );
  INVX1 U345 ( .A(n96), .Y(n295) );
  INVX1 U346 ( .A(n297), .Y(n296) );
  BUFX2 U347 ( .A(n433), .Y(n297) );
  AND2X2 U348 ( .A(n88), .B(n156), .Y(n298) );
  AND2X2 U349 ( .A(n164), .B(n138), .Y(n299) );
  INVX1 U350 ( .A(n299), .Y(n300) );
  AND2X1 U351 ( .A(n355), .B(n425), .Y(n301) );
  INVX1 U352 ( .A(n301), .Y(n302) );
  OR2X1 U353 ( .A(n315), .B(n442), .Y(n303) );
  INVX1 U354 ( .A(n304), .Y(n305) );
  AND2X2 U355 ( .A(n51), .B(n413), .Y(n306) );
  INVX1 U356 ( .A(n306), .Y(n307) );
  AND2X2 U357 ( .A(n431), .B(n28), .Y(n308) );
  INVX1 U358 ( .A(n40), .Y(n309) );
  AND2X2 U359 ( .A(n124), .B(n152), .Y(n312) );
  AND2X2 U360 ( .A(n81), .B(n128), .Y(n313) );
  AND2X2 U361 ( .A(n162), .B(n179), .Y(n314) );
  INVX1 U362 ( .A(n314), .Y(n315) );
  AND2X2 U363 ( .A(n355), .B(n175), .Y(n316) );
  INVX1 U364 ( .A(n316), .Y(n317) );
  INVX1 U365 ( .A(\Op<0> ), .Y(n352) );
  XNOR2X1 U366 ( .A(n328), .B(n341), .Y(n318) );
  INVX1 U367 ( .A(n318), .Y(n361) );
  INVX1 U368 ( .A(n7), .Y(n319) );
  AND2X2 U369 ( .A(n442), .B(n106), .Y(n320) );
  INVX1 U370 ( .A(n320), .Y(n439) );
  INVX1 U371 ( .A(n67), .Y(n322) );
  INVX1 U372 ( .A(\A<1> ), .Y(n325) );
  INVX1 U373 ( .A(n325), .Y(n326) );
  INVX4 U374 ( .A(n350), .Y(n452) );
  AND2X2 U375 ( .A(n316), .B(\sumOut<8> ), .Y(n327) );
  INVX1 U376 ( .A(n327), .Y(n441) );
  INVX1 U377 ( .A(\A<2> ), .Y(n328) );
  BUFX2 U378 ( .A(\B<7> ), .Y(n329) );
  BUFX2 U379 ( .A(\B<11> ), .Y(n330) );
  INVX1 U380 ( .A(n46), .Y(n337) );
  INVX1 U381 ( .A(n332), .Y(n437) );
  AOI21X1 U382 ( .A(n334), .B(n303), .C(n55), .Y(n333) );
  INVX1 U383 ( .A(n281), .Y(n375) );
  INVX1 U384 ( .A(n55), .Y(n445) );
  INVX1 U385 ( .A(n331), .Y(n335) );
  INVX1 U386 ( .A(n338), .Y(n336) );
  OR2X2 U387 ( .A(n34), .B(n63), .Y(n338) );
  INVX8 U388 ( .A(n340), .Y(n346) );
  INVX4 U389 ( .A(\Op<2> ), .Y(n442) );
  INVX4 U390 ( .A(n260), .Y(n425) );
  BUFX4 U391 ( .A(invB), .Y(n339) );
  BUFX4 U392 ( .A(invB), .Y(n340) );
  BUFX4 U393 ( .A(invA), .Y(n341) );
  XNOR2X1 U394 ( .A(\B<4> ), .B(n346), .Y(n488) );
  XNOR2X1 U395 ( .A(\B<5> ), .B(n346), .Y(n487) );
  INVX2 U396 ( .A(n345), .Y(n486) );
  XNOR2X1 U397 ( .A(\B<8> ), .B(n346), .Y(n484) );
  XNOR2X1 U398 ( .A(\B<10> ), .B(n346), .Y(n483) );
  XNOR2X1 U399 ( .A(\B<12> ), .B(n339), .Y(n384) );
  INVX2 U400 ( .A(n384), .Y(n481) );
  XNOR2X1 U401 ( .A(\B<15> ), .B(n339), .Y(n432) );
  INVX2 U402 ( .A(n432), .Y(\opB<15> ) );
  XNOR2X1 U403 ( .A(\A<1> ), .B(n14), .Y(n478) );
  XNOR2X1 U404 ( .A(\A<4> ), .B(n14), .Y(n475) );
  XNOR2X1 U405 ( .A(\A<5> ), .B(n14), .Y(n474) );
  XNOR2X1 U406 ( .A(\A<6> ), .B(n14), .Y(n473) );
  XNOR2X1 U407 ( .A(\A<9> ), .B(n14), .Y(n471) );
  XNOR2X1 U408 ( .A(\A<11> ), .B(n14), .Y(n469) );
  XNOR2X1 U409 ( .A(\A<12> ), .B(n341), .Y(n383) );
  XNOR2X1 U410 ( .A(\A<13> ), .B(n341), .Y(n409) );
  XNOR2X1 U411 ( .A(\A<14> ), .B(n14), .Y(n466) );
  XNOR2X1 U412 ( .A(n326), .B(n341), .Y(n427) );
  INVX2 U413 ( .A(n427), .Y(n455) );
  XNOR2X1 U414 ( .A(\A<3> ), .B(n341), .Y(n348) );
  XNOR2X1 U415 ( .A(\A<5> ), .B(n341), .Y(n395) );
  INVX2 U416 ( .A(n395), .Y(n458) );
  XNOR2X1 U417 ( .A(\A<6> ), .B(n341), .Y(n349) );
  XNOR2X1 U418 ( .A(\A<7> ), .B(n341), .Y(n350) );
  XNOR2X1 U419 ( .A(\A<8> ), .B(n341), .Y(n351) );
  XNOR2X1 U420 ( .A(\A<9> ), .B(n341), .Y(n401) );
  XNOR2X1 U421 ( .A(\A<14> ), .B(n341), .Y(n371) );
  NAND3X1 U422 ( .A(\Op<1> ), .B(\Op<2> ), .C(n352), .Y(n422) );
  INVX2 U423 ( .A(\Op<1> ), .Y(n355) );
  OAI21X1 U424 ( .A(n142), .B(n450), .C(n344), .Y(n353) );
  MUX2X1 U425 ( .B(n342), .A(n425), .S(n486), .Y(n354) );
  AOI21X1 U426 ( .A(\shiftOut<6> ), .B(n442), .C(n211), .Y(n356) );
  OAI21X1 U427 ( .A(n142), .B(n452), .C(n344), .Y(n357) );
  MUX2X1 U428 ( .B(n342), .A(n425), .S(n10), .Y(n358) );
  AOI21X1 U429 ( .A(\shiftOut<7> ), .B(n442), .C(n213), .Y(n359) );
  MUX2X1 U430 ( .B(n342), .A(n425), .S(n7), .Y(n360) );
  AOI21X1 U431 ( .A(n344), .B(n360), .C(n361), .Y(n365) );
  AOI21X1 U432 ( .A(n302), .B(n216), .C(n319), .Y(n364) );
  AND2X2 U433 ( .A(\sumOut<2> ), .B(n316), .Y(n363) );
  NOR3X1 U434 ( .A(n250), .B(n253), .C(n363), .Y(n366) );
  OAI21X1 U435 ( .A(n142), .B(n323), .C(n344), .Y(n367) );
  MUX2X1 U436 ( .B(n342), .A(n425), .S(n11), .Y(n368) );
  XNOR2X1 U437 ( .A(\B<14> ), .B(n340), .Y(n372) );
  INVX2 U438 ( .A(n372), .Y(n369) );
  MUX2X1 U439 ( .B(n342), .A(n425), .S(n369), .Y(n370) );
  AOI21X1 U440 ( .A(n302), .B(n220), .C(n372), .Y(n373) );
  AOI21X1 U441 ( .A(n446), .B(n218), .C(n202), .Y(n374) );
  OAI21X1 U442 ( .A(n375), .B(\sumOut<14> ), .C(n3), .Y(n376) );
  AND2X2 U443 ( .A(\sumOut<0> ), .B(n316), .Y(n381) );
  AOI21X1 U444 ( .A(n344), .B(n222), .C(n322), .Y(n380) );
  MUX2X1 U445 ( .B(n342), .A(n425), .S(n67), .Y(n378) );
  AOI21X1 U446 ( .A(n302), .B(n378), .C(n19), .Y(n379) );
  NOR3X1 U447 ( .A(n381), .B(n255), .C(n257), .Y(n438) );
  MUX2X1 U448 ( .B(n342), .A(n425), .S(n481), .Y(n382) );
  AOI21X1 U449 ( .A(n302), .B(n226), .C(n384), .Y(n385) );
  AOI21X1 U450 ( .A(n20), .B(n224), .C(n203), .Y(n386) );
  XNOR2X1 U451 ( .A(\B<10> ), .B(n340), .Y(n390) );
  INVX2 U452 ( .A(n390), .Y(n387) );
  MUX2X1 U453 ( .B(n342), .A(n425), .S(n387), .Y(n388) );
  AOI21X1 U454 ( .A(n302), .B(n230), .C(n390), .Y(n391) );
  AOI21X1 U455 ( .A(n449), .B(n228), .C(n204), .Y(n392) );
  AND2X2 U456 ( .A(n123), .B(n144), .Y(n393) );
  AND2X2 U457 ( .A(\shiftOut<5> ), .B(n442), .Y(n399) );
  XNOR2X1 U458 ( .A(n135), .B(n340), .Y(n394) );
  AOI21X1 U459 ( .A(n302), .B(n232), .C(n394), .Y(n398) );
  MUX2X1 U460 ( .B(n425), .A(n342), .S(n394), .Y(n396) );
  AOI21X1 U461 ( .A(n344), .B(n396), .C(n395), .Y(n397) );
  NOR3X1 U462 ( .A(n251), .B(n256), .C(n399), .Y(n440) );
  MUX2X1 U463 ( .B(n342), .A(n425), .S(n64), .Y(n400) );
  AOI21X1 U464 ( .A(n302), .B(n236), .C(n402), .Y(n403) );
  AOI21X1 U465 ( .A(n457), .B(n234), .C(n205), .Y(n404) );
  MUX2X1 U466 ( .B(n342), .A(n425), .S(\opB<15> ), .Y(n405) );
  OAI21X1 U467 ( .A(n142), .B(n13), .C(n344), .Y(n406) );
  AOI21X1 U468 ( .A(n13), .B(n238), .C(n407), .Y(n433) );
  MUX2X1 U469 ( .B(n342), .A(n425), .S(n15), .Y(n408) );
  AOI21X1 U470 ( .A(n302), .B(n242), .C(n410), .Y(n411) );
  AOI21X1 U471 ( .A(n467), .B(n240), .C(n206), .Y(n412) );
  OAI21X1 U472 ( .A(\sumOut<13> ), .B(n24), .C(n130), .Y(n413) );
  XNOR2X1 U473 ( .A(\B<4> ), .B(n340), .Y(n417) );
  INVX2 U474 ( .A(n417), .Y(n414) );
  MUX2X1 U475 ( .B(n342), .A(n425), .S(n414), .Y(n415) );
  AOI21X1 U476 ( .A(n302), .B(n246), .C(n417), .Y(n418) );
  AOI21X1 U477 ( .A(n39), .B(n244), .C(n207), .Y(n419) );
  OAI21X1 U478 ( .A(n142), .B(n451), .C(n344), .Y(n420) );
  MUX2X1 U479 ( .B(n342), .A(n425), .S(n456), .Y(n421) );
  OAI21X1 U480 ( .A(n142), .B(n35), .C(n302), .Y(n423) );
  MUX2X1 U481 ( .B(n342), .A(n425), .S(n12), .Y(n424) );
  MUX2X1 U482 ( .B(n342), .A(n425), .S(n60), .Y(n426) );
  AOI21X1 U483 ( .A(n302), .B(n248), .C(n59), .Y(n429) );
  AOI21X1 U484 ( .A(n455), .B(n95), .C(n209), .Y(n430) );
  NOR3X1 U485 ( .A(n97), .B(n287), .C(n258), .Y(n431) );
  NAND3X1 U486 ( .A(n332), .B(n308), .C(n306), .Y(n434) );
  NAND3X1 U487 ( .A(n70), .B(n432), .C(\sumOut<15> ), .Y(n436) );
  XNOR2X1 U488 ( .A(n262), .B(n46), .Y(N) );
  NOR3X1 U489 ( .A(n437), .B(n307), .C(n309), .Y(Z) );
  NAND3X1 U490 ( .A(n292), .B(n439), .C(n293), .Y(n462) );
  NAND3X1 U491 ( .A(n305), .B(n299), .C(n441), .Y(n447) );
  AOI21X1 U492 ( .A(n442), .B(n16), .C(n315), .Y(n443) );
endmodule


module alu_control ( .alu_op({\alu_op<2> , \alu_op<1> , \alu_op<0> }), inv_a, 
        inv_b, cin, .shamt({\shamt<3> , \shamt<2> , \shamt<1> , \shamt<0> }), 
        flip_1, flip_2, shift, SLBI, .opcode({\opcode<4> , \opcode<3> , 
        \opcode<2> , \opcode<1> , \opcode<0> }), .func({\func<1> , \func<0> }), 
    .immd({\immd<3> , \immd<2> , \immd<1> , \immd<0> }) );
  input \opcode<4> , \opcode<3> , \opcode<2> , \opcode<1> , \opcode<0> ,
         \func<1> , \func<0> , \immd<3> , \immd<2> , \immd<1> , \immd<0> ;
  output \alu_op<2> , \alu_op<1> , \alu_op<0> , inv_a, inv_b, cin, \shamt<3> ,
         \shamt<2> , \shamt<1> , \shamt<0> , flip_1, flip_2, shift, SLBI;
  wire   n97, n98, n1, n2, n3, n4, n5, n6, n7, n8, n9, n11, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n60,
         n61, n62, n63, n64, n65, n66, n67, n69, n71, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96;

  INVX1 U3 ( .A(\func<0> ), .Y(n76) );
  INVX1 U4 ( .A(n90), .Y(flip_1) );
  INVX1 U5 ( .A(\opcode<3> ), .Y(n1) );
  INVX1 U6 ( .A(n1), .Y(n2) );
  BUFX2 U7 ( .A(\opcode<1> ), .Y(n3) );
  BUFX2 U8 ( .A(n14), .Y(n4) );
  INVX1 U9 ( .A(\opcode<1> ), .Y(n5) );
  AND2X2 U10 ( .A(\opcode<4> ), .B(n74), .Y(n6) );
  INVX1 U11 ( .A(n4), .Y(n7) );
  INVX1 U12 ( .A(n85), .Y(n8) );
  INVX4 U13 ( .A(\opcode<2> ), .Y(n93) );
  INVX1 U14 ( .A(n14), .Y(n9) );
  INVX1 U15 ( .A(n14), .Y(n60) );
  AND2X2 U16 ( .A(\opcode<4> ), .B(n2), .Y(n55) );
  OR2X2 U17 ( .A(n36), .B(n11), .Y(shift) );
  OR2X2 U18 ( .A(n35), .B(n17), .Y(n11) );
  OR2X2 U19 ( .A(n65), .B(n13), .Y(\alu_op<2> ) );
  OR2X2 U20 ( .A(n63), .B(n64), .Y(n13) );
  OR2X2 U21 ( .A(n5), .B(\opcode<0> ), .Y(n14) );
  AND2X2 U22 ( .A(\opcode<4> ), .B(n74), .Y(n15) );
  INVX1 U23 ( .A(n6), .Y(n16) );
  AND2X2 U24 ( .A(n9), .B(n78), .Y(n17) );
  AND2X2 U25 ( .A(n78), .B(n7), .Y(n18) );
  INVX1 U26 ( .A(n18), .Y(n19) );
  AND2X2 U27 ( .A(n3), .B(\opcode<0> ), .Y(n20) );
  OR2X2 U28 ( .A(n62), .B(n85), .Y(n21) );
  INVX1 U29 ( .A(n21), .Y(n22) );
  AND2X2 U30 ( .A(n38), .B(n54), .Y(n23) );
  INVX1 U31 ( .A(n23), .Y(n24) );
  BUFX2 U32 ( .A(n84), .Y(n25) );
  AND2X2 U33 ( .A(\immd<3> ), .B(n34), .Y(n26) );
  INVX1 U34 ( .A(n26), .Y(n27) );
  AND2X2 U35 ( .A(n71), .B(n27), .Y(n28) );
  INVX1 U36 ( .A(n28), .Y(\shamt<3> ) );
  BUFX2 U37 ( .A(n87), .Y(n30) );
  AND2X2 U38 ( .A(n66), .B(n19), .Y(n31) );
  INVX1 U39 ( .A(n31), .Y(n32) );
  INVX1 U40 ( .A(n31), .Y(n33) );
  INVX1 U41 ( .A(n31), .Y(n34) );
  INVX1 U42 ( .A(n30), .Y(n35) );
  INVX1 U43 ( .A(n66), .Y(n36) );
  AND2X2 U44 ( .A(\opcode<2> ), .B(n6), .Y(n37) );
  AND2X2 U45 ( .A(n78), .B(n20), .Y(n38) );
  INVX1 U46 ( .A(flip_2), .Y(n90) );
  INVX1 U47 ( .A(\opcode<3> ), .Y(n74) );
  INVX1 U48 ( .A(n83), .Y(n39) );
  INVX1 U49 ( .A(n39), .Y(n40) );
  INVX1 U50 ( .A(n77), .Y(n41) );
  INVX1 U51 ( .A(n41), .Y(n42) );
  OR2X1 U52 ( .A(n66), .B(n85), .Y(n43) );
  INVX1 U53 ( .A(n43), .Y(n44) );
  OR2X1 U54 ( .A(n62), .B(n91), .Y(n45) );
  INVX1 U55 ( .A(n45), .Y(n46) );
  INVX1 U56 ( .A(n75), .Y(n78) );
  BUFX2 U57 ( .A(n86), .Y(n47) );
  BUFX2 U58 ( .A(n88), .Y(n48) );
  OR2X2 U59 ( .A(n53), .B(n19), .Y(n49) );
  INVX1 U60 ( .A(n49), .Y(n50) );
  OR2X1 U61 ( .A(n57), .B(n66), .Y(n51) );
  INVX1 U62 ( .A(n51), .Y(n52) );
  INVX1 U63 ( .A(n16), .Y(n92) );
  INVX1 U64 ( .A(n54), .Y(n53) );
  AND2X1 U65 ( .A(\func<0> ), .B(\func<1> ), .Y(n54) );
  INVX1 U66 ( .A(n55), .Y(n56) );
  INVX1 U67 ( .A(n20), .Y(n57) );
  AND2X2 U68 ( .A(n25), .B(n40), .Y(n58) );
  INVX1 U69 ( .A(n58), .Y(inv_a) );
  INVX1 U70 ( .A(n94), .Y(n61) );
  INVX1 U71 ( .A(n61), .Y(n62) );
  INVX1 U72 ( .A(n62), .Y(n63) );
  INVX1 U73 ( .A(n95), .Y(n64) );
  INVX1 U74 ( .A(n96), .Y(n65) );
  INVX1 U75 ( .A(n37), .Y(n66) );
  INVX1 U76 ( .A(n98), .Y(n67) );
  INVX1 U77 ( .A(n67), .Y(\alu_op<0> ) );
  INVX1 U78 ( .A(n97), .Y(n69) );
  INVX2 U79 ( .A(n69), .Y(\alu_op<1> ) );
  BUFX2 U80 ( .A(n30), .Y(n71) );
  INVX1 U81 ( .A(\opcode<4> ), .Y(n80) );
  BUFX2 U82 ( .A(inv_a), .Y(cin) );
  INVX1 U83 ( .A(n9), .Y(n91) );
  INVX1 U84 ( .A(\opcode<0> ), .Y(n85) );
  INVX1 U85 ( .A(n3), .Y(n82) );
  INVX1 U86 ( .A(n71), .Y(SLBI) );
  NAND3X1 U87 ( .A(n93), .B(n15), .C(n60), .Y(n87) );
  NAND3X1 U88 ( .A(\opcode<4> ), .B(\opcode<3> ), .C(n93), .Y(n75) );
  NAND3X1 U89 ( .A(\func<1> ), .B(n18), .C(n76), .Y(n77) );
  OAI21X1 U90 ( .A(n66), .B(n91), .C(n42), .Y(flip_2) );
  AND2X2 U91 ( .A(n33), .B(\immd<0> ), .Y(\shamt<0> ) );
  AND2X2 U92 ( .A(n32), .B(\immd<1> ), .Y(\shamt<1> ) );
  AND2X2 U93 ( .A(\immd<2> ), .B(n33), .Y(\shamt<2> ) );
  INVX2 U94 ( .A(\func<1> ), .Y(n79) );
  NAND3X1 U95 ( .A(\func<0> ), .B(n38), .C(n79), .Y(n84) );
  NAND3X1 U96 ( .A(n93), .B(n2), .C(n80), .Y(n94) );
  NOR3X1 U97 ( .A(n56), .B(n20), .C(n93), .Y(n81) );
  AOI21X1 U98 ( .A(n82), .B(n22), .C(n81), .Y(n83) );
  OAI21X1 U99 ( .A(n62), .B(n57), .C(n24), .Y(inv_b) );
  NOR3X1 U100 ( .A(inv_b), .B(n50), .C(n52), .Y(n89) );
  AOI21X1 U101 ( .A(\func<0> ), .B(n18), .C(n44), .Y(n86) );
  NAND3X1 U102 ( .A(n71), .B(n89), .C(n47), .Y(n98) );
  AOI21X1 U103 ( .A(\func<1> ), .B(n38), .C(n46), .Y(n88) );
  NAND3X1 U104 ( .A(n90), .B(n89), .C(n48), .Y(n97) );
  OAI21X1 U105 ( .A(n8), .B(\opcode<2> ), .C(n55), .Y(n96) );
  NAND3X1 U106 ( .A(n93), .B(n92), .C(n91), .Y(n95) );
endmodule


module reg3_5 ( .read({\read<2> , \read<1> , \read<0> }), .write({\write<2> , 
        \write<1> , \write<0> }), wr_en, rst, clk );
  input \write<2> , \write<1> , \write<0> , wr_en, rst, clk;
  output \read<2> , \read<1> , \read<0> ;
  wire   n1, n5, n9, n10, n11, n12, n13, n14, n15, n16;

  dff_451 d0 ( .q(\read<0> ), .d(n16), .clk(clk), .rst(rst) );
  dff_450 d1 ( .q(\read<1> ), .d(n15), .clk(clk), .rst(rst) );
  dff_449 d2 ( .q(\read<2> ), .d(n14), .clk(clk), .rst(rst) );
  AOI22X1 U5 ( .A(\read<2> ), .B(n10), .C(\write<2> ), .D(wr_en), .Y(n13) );
  AOI22X1 U6 ( .A(\read<1> ), .B(n10), .C(\write<1> ), .D(wr_en), .Y(n12) );
  AOI22X1 U7 ( .A(\read<0> ), .B(n10), .C(\write<0> ), .D(wr_en), .Y(n11) );
  INVX1 U1 ( .A(wr_en), .Y(n10) );
  BUFX2 U2 ( .A(n11), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(n16) );
  BUFX2 U4 ( .A(n12), .Y(n5) );
  INVX1 U8 ( .A(n5), .Y(n15) );
  BUFX2 U9 ( .A(n13), .Y(n9) );
  INVX1 U10 ( .A(n9), .Y(n14) );
endmodule


module reg3_4 ( .read({\read<2> , \read<1> , \read<0> }), .write({\write<2> , 
        \write<1> , \write<0> }), wr_en, rst, clk );
  input \write<2> , \write<1> , \write<0> , wr_en, rst, clk;
  output \read<2> , \read<1> , \read<0> ;
  wire   n1, n5, n9, n10, n11, n12, n13, n14, n15, n16;

  dff_448 d0 ( .q(\read<0> ), .d(n16), .clk(clk), .rst(rst) );
  dff_447 d1 ( .q(\read<1> ), .d(n15), .clk(clk), .rst(rst) );
  dff_446 d2 ( .q(\read<2> ), .d(n14), .clk(clk), .rst(rst) );
  AOI22X1 U5 ( .A(\read<2> ), .B(n10), .C(\write<2> ), .D(wr_en), .Y(n13) );
  AOI22X1 U6 ( .A(\read<1> ), .B(n10), .C(\write<1> ), .D(wr_en), .Y(n12) );
  AOI22X1 U7 ( .A(\read<0> ), .B(n10), .C(\write<0> ), .D(wr_en), .Y(n11) );
  INVX1 U1 ( .A(wr_en), .Y(n10) );
  BUFX2 U2 ( .A(n11), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(n16) );
  BUFX2 U4 ( .A(n12), .Y(n5) );
  INVX1 U8 ( .A(n5), .Y(n15) );
  BUFX2 U9 ( .A(n13), .Y(n9) );
  INVX1 U10 ( .A(n9), .Y(n14) );
endmodule


module reg3_3 ( .read({\read<2> , \read<1> , \read<0> }), .write({\write<2> , 
        \write<1> , \write<0> }), wr_en, rst, clk );
  input \write<2> , \write<1> , \write<0> , wr_en, rst, clk;
  output \read<2> , \read<1> , \read<0> ;
  wire   n1, n5, n9, n10, n11, n12, n13, n14, n15, n16;

  dff_445 d0 ( .q(\read<0> ), .d(n16), .clk(clk), .rst(rst) );
  dff_444 d1 ( .q(\read<1> ), .d(n15), .clk(clk), .rst(rst) );
  dff_443 d2 ( .q(\read<2> ), .d(n14), .clk(clk), .rst(rst) );
  AOI22X1 U5 ( .A(\read<2> ), .B(n10), .C(\write<2> ), .D(wr_en), .Y(n13) );
  AOI22X1 U6 ( .A(\read<1> ), .B(n10), .C(\write<1> ), .D(wr_en), .Y(n12) );
  AOI22X1 U7 ( .A(\read<0> ), .B(n10), .C(\write<0> ), .D(wr_en), .Y(n11) );
  INVX1 U1 ( .A(wr_en), .Y(n10) );
  BUFX2 U2 ( .A(n11), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(n16) );
  BUFX2 U4 ( .A(n12), .Y(n5) );
  INVX1 U8 ( .A(n5), .Y(n15) );
  BUFX2 U9 ( .A(n13), .Y(n9) );
  INVX1 U10 ( .A(n9), .Y(n14) );
endmodule


module reg16_25 ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n1, n18, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91;

  dff_442 d0 ( .q(\read<0> ), .d(n91), .clk(clk), .rst(rst) );
  dff_441 d1 ( .q(\read<1> ), .d(n90), .clk(clk), .rst(rst) );
  dff_440 d2 ( .q(\read<2> ), .d(n89), .clk(clk), .rst(rst) );
  dff_439 d3 ( .q(\read<3> ), .d(n88), .clk(clk), .rst(rst) );
  dff_438 d4 ( .q(\read<4> ), .d(n87), .clk(clk), .rst(rst) );
  dff_437 d5 ( .q(\read<5> ), .d(n86), .clk(clk), .rst(rst) );
  dff_436 d6 ( .q(\read<6> ), .d(n85), .clk(clk), .rst(rst) );
  dff_435 d7 ( .q(\read<7> ), .d(n84), .clk(clk), .rst(rst) );
  dff_434 d8 ( .q(\read<8> ), .d(n83), .clk(clk), .rst(rst) );
  dff_433 d9 ( .q(\read<9> ), .d(n82), .clk(clk), .rst(rst) );
  dff_432 d10 ( .q(\read<10> ), .d(n81), .clk(clk), .rst(rst) );
  dff_431 d11 ( .q(\read<11> ), .d(n80), .clk(clk), .rst(rst) );
  dff_430 d12 ( .q(\read<12> ), .d(n79), .clk(clk), .rst(rst) );
  dff_429 d13 ( .q(\read<13> ), .d(n78), .clk(clk), .rst(rst) );
  dff_428 d14 ( .q(\read<14> ), .d(n77), .clk(clk), .rst(rst) );
  dff_427 d15 ( .q(\read<15> ), .d(n76), .clk(clk), .rst(rst) );
  AOI22X1 U18 ( .A(\read<9> ), .B(n58), .C(\write<9> ), .D(n56), .Y(n75) );
  AOI22X1 U19 ( .A(\read<8> ), .B(n58), .C(\write<8> ), .D(n56), .Y(n74) );
  AOI22X1 U20 ( .A(\read<7> ), .B(n58), .C(\write<7> ), .D(n56), .Y(n73) );
  AOI22X1 U21 ( .A(\read<6> ), .B(n58), .C(\write<6> ), .D(n56), .Y(n72) );
  AOI22X1 U22 ( .A(\read<5> ), .B(n59), .C(\write<5> ), .D(n56), .Y(n71) );
  AOI22X1 U23 ( .A(\read<4> ), .B(n59), .C(\write<4> ), .D(n56), .Y(n70) );
  AOI22X1 U24 ( .A(\read<3> ), .B(n59), .C(\write<3> ), .D(n56), .Y(n69) );
  AOI22X1 U25 ( .A(\read<2> ), .B(n59), .C(\write<2> ), .D(n56), .Y(n68) );
  AOI22X1 U26 ( .A(\read<1> ), .B(n59), .C(\write<1> ), .D(n56), .Y(n67) );
  AOI22X1 U27 ( .A(n50), .B(n59), .C(\write<15> ), .D(n56), .Y(n66) );
  AOI22X1 U28 ( .A(n49), .B(n59), .C(\write<14> ), .D(n56), .Y(n65) );
  AOI22X1 U29 ( .A(n51), .B(n59), .C(\write<13> ), .D(n56), .Y(n64) );
  AOI22X1 U30 ( .A(n53), .B(n59), .C(\write<12> ), .D(n57), .Y(n63) );
  AOI22X1 U31 ( .A(n52), .B(n59), .C(\write<11> ), .D(n57), .Y(n62) );
  AOI22X1 U32 ( .A(\read<10> ), .B(n59), .C(\write<10> ), .D(n57), .Y(n61) );
  AOI22X1 U33 ( .A(\read<0> ), .B(n59), .C(\write<0> ), .D(n57), .Y(n60) );
  INVX1 U1 ( .A(wr_en), .Y(n55) );
  INVX1 U2 ( .A(n54), .Y(n58) );
  INVX1 U3 ( .A(n55), .Y(n54) );
  INVX1 U4 ( .A(n58), .Y(n57) );
  INVX1 U5 ( .A(n54), .Y(n59) );
  INVX1 U6 ( .A(n58), .Y(n56) );
  BUFX2 U7 ( .A(n60), .Y(n1) );
  INVX1 U8 ( .A(n1), .Y(n91) );
  BUFX2 U9 ( .A(n61), .Y(n18) );
  INVX1 U10 ( .A(n18), .Y(n81) );
  BUFX2 U11 ( .A(n62), .Y(n35) );
  INVX1 U12 ( .A(n35), .Y(n80) );
  BUFX2 U13 ( .A(n63), .Y(n36) );
  INVX1 U14 ( .A(n36), .Y(n79) );
  BUFX2 U15 ( .A(n64), .Y(n37) );
  INVX1 U16 ( .A(n37), .Y(n78) );
  BUFX2 U17 ( .A(n65), .Y(n38) );
  INVX1 U34 ( .A(n38), .Y(n77) );
  BUFX2 U35 ( .A(n66), .Y(n39) );
  INVX1 U36 ( .A(n39), .Y(n76) );
  BUFX2 U37 ( .A(n67), .Y(n40) );
  INVX1 U38 ( .A(n40), .Y(n90) );
  BUFX2 U39 ( .A(n68), .Y(n41) );
  INVX1 U40 ( .A(n41), .Y(n89) );
  BUFX2 U41 ( .A(n69), .Y(n42) );
  INVX1 U42 ( .A(n42), .Y(n88) );
  BUFX2 U43 ( .A(n70), .Y(n43) );
  INVX1 U44 ( .A(n43), .Y(n87) );
  BUFX2 U45 ( .A(n71), .Y(n44) );
  INVX1 U46 ( .A(n44), .Y(n86) );
  BUFX2 U47 ( .A(n72), .Y(n45) );
  INVX1 U48 ( .A(n45), .Y(n85) );
  BUFX2 U49 ( .A(n73), .Y(n46) );
  INVX1 U50 ( .A(n46), .Y(n84) );
  BUFX2 U51 ( .A(n74), .Y(n47) );
  INVX1 U52 ( .A(n47), .Y(n83) );
  BUFX2 U53 ( .A(n75), .Y(n48) );
  INVX1 U54 ( .A(n48), .Y(n82) );
  BUFX2 U55 ( .A(\read<14> ), .Y(n49) );
  BUFX2 U56 ( .A(\read<15> ), .Y(n50) );
  BUFX2 U57 ( .A(\read<13> ), .Y(n51) );
  BUFX2 U58 ( .A(\read<11> ), .Y(n52) );
  BUFX2 U59 ( .A(\read<12> ), .Y(n53) );
endmodule


module reg16_24 ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52;

  dff_426 d0 ( .q(\read<0> ), .d(n37), .clk(clk), .rst(rst) );
  dff_425 d1 ( .q(\read<1> ), .d(n38), .clk(clk), .rst(rst) );
  dff_424 d2 ( .q(\read<2> ), .d(n39), .clk(clk), .rst(rst) );
  dff_423 d3 ( .q(\read<3> ), .d(n40), .clk(clk), .rst(rst) );
  dff_422 d4 ( .q(\read<4> ), .d(n41), .clk(clk), .rst(rst) );
  dff_421 d5 ( .q(\read<5> ), .d(n42), .clk(clk), .rst(rst) );
  dff_420 d6 ( .q(\read<6> ), .d(n43), .clk(clk), .rst(rst) );
  dff_419 d7 ( .q(\read<7> ), .d(n44), .clk(clk), .rst(rst) );
  dff_418 d8 ( .q(\read<8> ), .d(n45), .clk(clk), .rst(rst) );
  dff_417 d9 ( .q(\read<9> ), .d(n46), .clk(clk), .rst(rst) );
  dff_416 d10 ( .q(\read<10> ), .d(n47), .clk(clk), .rst(rst) );
  dff_415 d11 ( .q(\read<11> ), .d(n48), .clk(clk), .rst(rst) );
  dff_414 d12 ( .q(\read<12> ), .d(n49), .clk(clk), .rst(rst) );
  dff_413 d13 ( .q(\read<13> ), .d(n50), .clk(clk), .rst(rst) );
  dff_412 d14 ( .q(\read<14> ), .d(n51), .clk(clk), .rst(rst) );
  dff_411 d15 ( .q(\read<15> ), .d(n52), .clk(clk), .rst(rst) );
  INVX1 U1 ( .A(\write<4> ), .Y(n27) );
  INVX1 U2 ( .A(\read<4> ), .Y(n28) );
  INVX1 U3 ( .A(\read<5> ), .Y(n26) );
  INVX1 U4 ( .A(\read<6> ), .Y(n24) );
  INVX1 U5 ( .A(\read<7> ), .Y(n22) );
  INVX1 U6 ( .A(\read<8> ), .Y(n20) );
  INVX1 U7 ( .A(\read<9> ), .Y(n18) );
  INVX1 U8 ( .A(\read<10> ), .Y(n16) );
  INVX1 U9 ( .A(\read<11> ), .Y(n14) );
  INVX1 U10 ( .A(\write<12> ), .Y(n11) );
  INVX1 U11 ( .A(\read<12> ), .Y(n12) );
  INVX1 U12 ( .A(\write<13> ), .Y(n9) );
  INVX1 U13 ( .A(\read<13> ), .Y(n10) );
  INVX1 U14 ( .A(\read<14> ), .Y(n8) );
  INVX1 U15 ( .A(\read<15> ), .Y(n6) );
  INVX1 U16 ( .A(\read<0> ), .Y(n36) );
  INVX1 U17 ( .A(\read<1> ), .Y(n34) );
  INVX1 U18 ( .A(\read<2> ), .Y(n32) );
  INVX1 U19 ( .A(\read<3> ), .Y(n30) );
  INVX1 U20 ( .A(n4), .Y(n2) );
  INVX1 U21 ( .A(wr_en), .Y(n4) );
  INVX1 U22 ( .A(n4), .Y(n3) );
  INVX1 U23 ( .A(n3), .Y(n1) );
  INVX1 U24 ( .A(\write<1> ), .Y(n33) );
  INVX1 U25 ( .A(\write<0> ), .Y(n35) );
  MUX2X1 U26 ( .B(n26), .A(n25), .S(n2), .Y(n42) );
  INVX1 U27 ( .A(\write<8> ), .Y(n19) );
  MUX2X1 U28 ( .B(n21), .A(n22), .S(n4), .Y(n44) );
  INVX1 U29 ( .A(\write<3> ), .Y(n29) );
  INVX1 U30 ( .A(\write<6> ), .Y(n23) );
  MUX2X1 U31 ( .B(n5), .A(n6), .S(n1), .Y(n52) );
  MUX2X1 U32 ( .B(n7), .A(n8), .S(n1), .Y(n51) );
  INVX1 U33 ( .A(\write<2> ), .Y(n31) );
  INVX1 U34 ( .A(\write<5> ), .Y(n25) );
  INVX1 U35 ( .A(\write<14> ), .Y(n7) );
  INVX1 U36 ( .A(\write<11> ), .Y(n13) );
  INVX1 U37 ( .A(\write<10> ), .Y(n15) );
  INVX1 U38 ( .A(\write<9> ), .Y(n17) );
  INVX1 U39 ( .A(\write<15> ), .Y(n5) );
  INVX1 U40 ( .A(\write<7> ), .Y(n21) );
  MUX2X1 U41 ( .B(n10), .A(n9), .S(n3), .Y(n50) );
  MUX2X1 U42 ( .B(n12), .A(n11), .S(n3), .Y(n49) );
  MUX2X1 U43 ( .B(n14), .A(n13), .S(n2), .Y(n48) );
  MUX2X1 U44 ( .B(n16), .A(n15), .S(n2), .Y(n47) );
  MUX2X1 U45 ( .B(n18), .A(n17), .S(n2), .Y(n46) );
  MUX2X1 U46 ( .B(n20), .A(n19), .S(n2), .Y(n45) );
  MUX2X1 U47 ( .B(n24), .A(n23), .S(n2), .Y(n43) );
  MUX2X1 U48 ( .B(n28), .A(n27), .S(n2), .Y(n41) );
  MUX2X1 U49 ( .B(n30), .A(n29), .S(n2), .Y(n40) );
  MUX2X1 U50 ( .B(n32), .A(n31), .S(n2), .Y(n39) );
  MUX2X1 U51 ( .B(n34), .A(n33), .S(n2), .Y(n38) );
  MUX2X1 U52 ( .B(n36), .A(n35), .S(n2), .Y(n37) );
endmodule


module reg16_23 ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n1, n18, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86;

  dff_410 d0 ( .q(\read<0> ), .d(n86), .clk(clk), .rst(rst) );
  dff_409 d1 ( .q(\read<1> ), .d(n85), .clk(clk), .rst(rst) );
  dff_408 d2 ( .q(\read<2> ), .d(n84), .clk(clk), .rst(rst) );
  dff_407 d3 ( .q(\read<3> ), .d(n83), .clk(clk), .rst(rst) );
  dff_406 d4 ( .q(\read<4> ), .d(n82), .clk(clk), .rst(rst) );
  dff_405 d5 ( .q(\read<5> ), .d(n81), .clk(clk), .rst(rst) );
  dff_404 d6 ( .q(\read<6> ), .d(n80), .clk(clk), .rst(rst) );
  dff_403 d7 ( .q(\read<7> ), .d(n79), .clk(clk), .rst(rst) );
  dff_402 d8 ( .q(\read<8> ), .d(n78), .clk(clk), .rst(rst) );
  dff_401 d9 ( .q(\read<9> ), .d(n77), .clk(clk), .rst(rst) );
  dff_400 d10 ( .q(\read<10> ), .d(n76), .clk(clk), .rst(rst) );
  dff_399 d11 ( .q(\read<11> ), .d(n75), .clk(clk), .rst(rst) );
  dff_398 d12 ( .q(\read<12> ), .d(n74), .clk(clk), .rst(rst) );
  dff_397 d13 ( .q(\read<13> ), .d(n73), .clk(clk), .rst(rst) );
  dff_396 d14 ( .q(\read<14> ), .d(n72), .clk(clk), .rst(rst) );
  dff_395 d15 ( .q(\read<15> ), .d(n71), .clk(clk), .rst(rst) );
  AOI22X1 U18 ( .A(\read<9> ), .B(n53), .C(\write<9> ), .D(n51), .Y(n70) );
  AOI22X1 U19 ( .A(\read<8> ), .B(n53), .C(\write<8> ), .D(n51), .Y(n69) );
  AOI22X1 U20 ( .A(\read<7> ), .B(n53), .C(\write<7> ), .D(n51), .Y(n68) );
  AOI22X1 U21 ( .A(\read<6> ), .B(n53), .C(\write<6> ), .D(n51), .Y(n67) );
  AOI22X1 U22 ( .A(\read<5> ), .B(n54), .C(\write<5> ), .D(n51), .Y(n66) );
  AOI22X1 U23 ( .A(\read<4> ), .B(n54), .C(\write<4> ), .D(n51), .Y(n65) );
  AOI22X1 U24 ( .A(\read<3> ), .B(n54), .C(\write<3> ), .D(n51), .Y(n64) );
  AOI22X1 U25 ( .A(\read<2> ), .B(n54), .C(\write<2> ), .D(n51), .Y(n63) );
  AOI22X1 U26 ( .A(\read<1> ), .B(n54), .C(\write<1> ), .D(n51), .Y(n62) );
  AOI22X1 U27 ( .A(\read<15> ), .B(n54), .C(\write<15> ), .D(n51), .Y(n61) );
  AOI22X1 U28 ( .A(\read<14> ), .B(n54), .C(\write<14> ), .D(n51), .Y(n60) );
  AOI22X1 U29 ( .A(\read<13> ), .B(n54), .C(\write<13> ), .D(n51), .Y(n59) );
  AOI22X1 U30 ( .A(\read<12> ), .B(n54), .C(\write<12> ), .D(n52), .Y(n58) );
  AOI22X1 U31 ( .A(\read<11> ), .B(n54), .C(\write<11> ), .D(n52), .Y(n57) );
  AOI22X1 U32 ( .A(\read<10> ), .B(n54), .C(\write<10> ), .D(n52), .Y(n56) );
  AOI22X1 U33 ( .A(\read<0> ), .B(n54), .C(\write<0> ), .D(n52), .Y(n55) );
  INVX1 U1 ( .A(wr_en), .Y(n50) );
  INVX1 U2 ( .A(n49), .Y(n53) );
  INVX1 U3 ( .A(n50), .Y(n49) );
  INVX1 U4 ( .A(n49), .Y(n54) );
  INVX1 U5 ( .A(n53), .Y(n52) );
  INVX1 U6 ( .A(n53), .Y(n51) );
  BUFX2 U7 ( .A(n55), .Y(n1) );
  INVX1 U8 ( .A(n1), .Y(n86) );
  BUFX2 U9 ( .A(n56), .Y(n18) );
  INVX1 U10 ( .A(n18), .Y(n76) );
  BUFX2 U11 ( .A(n57), .Y(n35) );
  INVX1 U12 ( .A(n35), .Y(n75) );
  BUFX2 U13 ( .A(n58), .Y(n36) );
  INVX1 U14 ( .A(n36), .Y(n74) );
  BUFX2 U15 ( .A(n59), .Y(n37) );
  INVX1 U16 ( .A(n37), .Y(n73) );
  BUFX2 U17 ( .A(n60), .Y(n38) );
  INVX1 U34 ( .A(n38), .Y(n72) );
  BUFX2 U35 ( .A(n61), .Y(n39) );
  INVX1 U36 ( .A(n39), .Y(n71) );
  BUFX2 U37 ( .A(n62), .Y(n40) );
  INVX1 U38 ( .A(n40), .Y(n85) );
  BUFX2 U39 ( .A(n63), .Y(n41) );
  INVX1 U40 ( .A(n41), .Y(n84) );
  BUFX2 U41 ( .A(n64), .Y(n42) );
  INVX1 U42 ( .A(n42), .Y(n83) );
  BUFX2 U43 ( .A(n65), .Y(n43) );
  INVX1 U44 ( .A(n43), .Y(n82) );
  BUFX2 U45 ( .A(n66), .Y(n44) );
  INVX1 U46 ( .A(n44), .Y(n81) );
  BUFX2 U47 ( .A(n67), .Y(n45) );
  INVX1 U48 ( .A(n45), .Y(n80) );
  BUFX2 U49 ( .A(n68), .Y(n46) );
  INVX1 U50 ( .A(n46), .Y(n79) );
  BUFX2 U51 ( .A(n69), .Y(n47) );
  INVX1 U52 ( .A(n47), .Y(n78) );
  BUFX2 U53 ( .A(n70), .Y(n48) );
  INVX1 U54 ( .A(n48), .Y(n77) );
endmodule


module reg16_22 ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n1, n18, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84;

  dff_394 d0 ( .q(\read<0> ), .d(n84), .clk(clk), .rst(rst) );
  dff_393 d1 ( .q(\read<1> ), .d(n83), .clk(clk), .rst(rst) );
  dff_392 d2 ( .q(\read<2> ), .d(n82), .clk(clk), .rst(rst) );
  dff_391 d3 ( .q(\read<3> ), .d(n81), .clk(clk), .rst(rst) );
  dff_390 d4 ( .q(\read<4> ), .d(n80), .clk(clk), .rst(rst) );
  dff_389 d5 ( .q(\read<5> ), .d(n79), .clk(clk), .rst(rst) );
  dff_388 d6 ( .q(\read<6> ), .d(n78), .clk(clk), .rst(rst) );
  dff_387 d7 ( .q(\read<7> ), .d(n77), .clk(clk), .rst(rst) );
  dff_386 d8 ( .q(\read<8> ), .d(n76), .clk(clk), .rst(rst) );
  dff_385 d9 ( .q(\read<9> ), .d(n75), .clk(clk), .rst(rst) );
  dff_384 d10 ( .q(\read<10> ), .d(n74), .clk(clk), .rst(rst) );
  dff_383 d11 ( .q(\read<11> ), .d(n73), .clk(clk), .rst(rst) );
  dff_382 d12 ( .q(\read<12> ), .d(n72), .clk(clk), .rst(rst) );
  dff_381 d13 ( .q(\read<13> ), .d(n71), .clk(clk), .rst(rst) );
  dff_380 d14 ( .q(\read<14> ), .d(n70), .clk(clk), .rst(rst) );
  dff_379 d15 ( .q(\read<15> ), .d(n69), .clk(clk), .rst(rst) );
  AOI22X1 U18 ( .A(\read<9> ), .B(n49), .C(\write<9> ), .D(n50), .Y(n68) );
  AOI22X1 U19 ( .A(\read<8> ), .B(n49), .C(\write<8> ), .D(n50), .Y(n67) );
  AOI22X1 U20 ( .A(\read<7> ), .B(n49), .C(\write<7> ), .D(n50), .Y(n66) );
  AOI22X1 U21 ( .A(\read<6> ), .B(n49), .C(\write<6> ), .D(n50), .Y(n65) );
  AOI22X1 U22 ( .A(\read<5> ), .B(n52), .C(\write<5> ), .D(n50), .Y(n64) );
  AOI22X1 U23 ( .A(\read<4> ), .B(n52), .C(\write<4> ), .D(n50), .Y(n63) );
  AOI22X1 U24 ( .A(\read<3> ), .B(n52), .C(\write<3> ), .D(n50), .Y(n62) );
  AOI22X1 U25 ( .A(\read<2> ), .B(n52), .C(\write<2> ), .D(n50), .Y(n61) );
  AOI22X1 U26 ( .A(\read<1> ), .B(n52), .C(\write<1> ), .D(n50), .Y(n60) );
  AOI22X1 U27 ( .A(\read<15> ), .B(n52), .C(\write<15> ), .D(n50), .Y(n59) );
  AOI22X1 U28 ( .A(\read<14> ), .B(n52), .C(\write<14> ), .D(n50), .Y(n58) );
  AOI22X1 U29 ( .A(\read<13> ), .B(n52), .C(\write<13> ), .D(n50), .Y(n57) );
  AOI22X1 U30 ( .A(\read<12> ), .B(n52), .C(\write<12> ), .D(n51), .Y(n56) );
  AOI22X1 U31 ( .A(\read<11> ), .B(n52), .C(\write<11> ), .D(n51), .Y(n55) );
  AOI22X1 U32 ( .A(\read<10> ), .B(n52), .C(\write<10> ), .D(n51), .Y(n54) );
  AOI22X1 U33 ( .A(\read<0> ), .B(n52), .C(\write<0> ), .D(n51), .Y(n53) );
  INVX1 U1 ( .A(wr_en), .Y(n49) );
  INVX1 U2 ( .A(wr_en), .Y(n52) );
  INVX1 U3 ( .A(n49), .Y(n51) );
  INVX1 U4 ( .A(n49), .Y(n50) );
  BUFX2 U5 ( .A(n53), .Y(n1) );
  INVX1 U6 ( .A(n1), .Y(n84) );
  BUFX2 U7 ( .A(n54), .Y(n18) );
  INVX1 U8 ( .A(n18), .Y(n74) );
  BUFX2 U9 ( .A(n55), .Y(n35) );
  INVX1 U10 ( .A(n35), .Y(n73) );
  BUFX2 U11 ( .A(n56), .Y(n36) );
  INVX1 U12 ( .A(n36), .Y(n72) );
  BUFX2 U13 ( .A(n57), .Y(n37) );
  INVX1 U14 ( .A(n37), .Y(n71) );
  BUFX2 U15 ( .A(n58), .Y(n38) );
  INVX1 U16 ( .A(n38), .Y(n70) );
  BUFX2 U17 ( .A(n59), .Y(n39) );
  INVX1 U34 ( .A(n39), .Y(n69) );
  BUFX2 U35 ( .A(n60), .Y(n40) );
  INVX1 U36 ( .A(n40), .Y(n83) );
  BUFX2 U37 ( .A(n61), .Y(n41) );
  INVX1 U38 ( .A(n41), .Y(n82) );
  BUFX2 U39 ( .A(n62), .Y(n42) );
  INVX1 U40 ( .A(n42), .Y(n81) );
  BUFX2 U41 ( .A(n63), .Y(n43) );
  INVX1 U42 ( .A(n43), .Y(n80) );
  BUFX2 U43 ( .A(n64), .Y(n44) );
  INVX1 U44 ( .A(n44), .Y(n79) );
  BUFX2 U45 ( .A(n65), .Y(n45) );
  INVX1 U46 ( .A(n45), .Y(n78) );
  BUFX2 U47 ( .A(n66), .Y(n46) );
  INVX1 U48 ( .A(n46), .Y(n77) );
  BUFX2 U49 ( .A(n67), .Y(n47) );
  INVX1 U50 ( .A(n47), .Y(n76) );
  BUFX2 U51 ( .A(n68), .Y(n48) );
  INVX1 U52 ( .A(n48), .Y(n75) );
endmodule


module reg16_21 ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n1, n18, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84;

  dff_378 d0 ( .q(\read<0> ), .d(n84), .clk(clk), .rst(rst) );
  dff_377 d1 ( .q(\read<1> ), .d(n83), .clk(clk), .rst(rst) );
  dff_376 d2 ( .q(\read<2> ), .d(n82), .clk(clk), .rst(rst) );
  dff_375 d3 ( .q(\read<3> ), .d(n81), .clk(clk), .rst(rst) );
  dff_374 d4 ( .q(\read<4> ), .d(n80), .clk(clk), .rst(rst) );
  dff_373 d5 ( .q(\read<5> ), .d(n79), .clk(clk), .rst(rst) );
  dff_372 d6 ( .q(\read<6> ), .d(n78), .clk(clk), .rst(rst) );
  dff_371 d7 ( .q(\read<7> ), .d(n77), .clk(clk), .rst(rst) );
  dff_370 d8 ( .q(\read<8> ), .d(n76), .clk(clk), .rst(rst) );
  dff_369 d9 ( .q(\read<9> ), .d(n75), .clk(clk), .rst(rst) );
  dff_368 d10 ( .q(\read<10> ), .d(n74), .clk(clk), .rst(rst) );
  dff_367 d11 ( .q(\read<11> ), .d(n73), .clk(clk), .rst(rst) );
  dff_366 d12 ( .q(\read<12> ), .d(n72), .clk(clk), .rst(rst) );
  dff_365 d13 ( .q(\read<13> ), .d(n71), .clk(clk), .rst(rst) );
  dff_364 d14 ( .q(\read<14> ), .d(n70), .clk(clk), .rst(rst) );
  dff_363 d15 ( .q(\read<15> ), .d(n69), .clk(clk), .rst(rst) );
  AOI22X1 U18 ( .A(\read<9> ), .B(n49), .C(\write<9> ), .D(n50), .Y(n68) );
  AOI22X1 U19 ( .A(\read<8> ), .B(n49), .C(\write<8> ), .D(n50), .Y(n67) );
  AOI22X1 U20 ( .A(\read<7> ), .B(n49), .C(\write<7> ), .D(n50), .Y(n66) );
  AOI22X1 U21 ( .A(\read<6> ), .B(n49), .C(\write<6> ), .D(n50), .Y(n65) );
  AOI22X1 U22 ( .A(\read<5> ), .B(n52), .C(\write<5> ), .D(n50), .Y(n64) );
  AOI22X1 U23 ( .A(\read<4> ), .B(n52), .C(\write<4> ), .D(n50), .Y(n63) );
  AOI22X1 U24 ( .A(\read<3> ), .B(n52), .C(\write<3> ), .D(n50), .Y(n62) );
  AOI22X1 U25 ( .A(\read<2> ), .B(n52), .C(\write<2> ), .D(n50), .Y(n61) );
  AOI22X1 U26 ( .A(\read<1> ), .B(n52), .C(\write<1> ), .D(n50), .Y(n60) );
  AOI22X1 U27 ( .A(\read<15> ), .B(n52), .C(\write<15> ), .D(n50), .Y(n59) );
  AOI22X1 U28 ( .A(\read<14> ), .B(n52), .C(\write<14> ), .D(n50), .Y(n58) );
  AOI22X1 U29 ( .A(\read<13> ), .B(n52), .C(\write<13> ), .D(n50), .Y(n57) );
  AOI22X1 U30 ( .A(\read<12> ), .B(n52), .C(\write<12> ), .D(n51), .Y(n56) );
  AOI22X1 U31 ( .A(\read<11> ), .B(n52), .C(\write<11> ), .D(n51), .Y(n55) );
  AOI22X1 U32 ( .A(\read<10> ), .B(n52), .C(\write<10> ), .D(n51), .Y(n54) );
  AOI22X1 U33 ( .A(\read<0> ), .B(n52), .C(\write<0> ), .D(n51), .Y(n53) );
  INVX1 U1 ( .A(wr_en), .Y(n49) );
  INVX1 U2 ( .A(n49), .Y(n51) );
  INVX1 U3 ( .A(wr_en), .Y(n52) );
  INVX1 U4 ( .A(n49), .Y(n50) );
  BUFX2 U5 ( .A(n53), .Y(n1) );
  INVX1 U6 ( .A(n1), .Y(n84) );
  BUFX2 U7 ( .A(n54), .Y(n18) );
  INVX1 U8 ( .A(n18), .Y(n74) );
  BUFX2 U9 ( .A(n55), .Y(n35) );
  INVX1 U10 ( .A(n35), .Y(n73) );
  BUFX2 U11 ( .A(n56), .Y(n36) );
  INVX1 U12 ( .A(n36), .Y(n72) );
  BUFX2 U13 ( .A(n57), .Y(n37) );
  INVX1 U14 ( .A(n37), .Y(n71) );
  BUFX2 U15 ( .A(n58), .Y(n38) );
  INVX1 U16 ( .A(n38), .Y(n70) );
  BUFX2 U17 ( .A(n59), .Y(n39) );
  INVX1 U34 ( .A(n39), .Y(n69) );
  BUFX2 U35 ( .A(n60), .Y(n40) );
  INVX1 U36 ( .A(n40), .Y(n83) );
  BUFX2 U37 ( .A(n61), .Y(n41) );
  INVX1 U38 ( .A(n41), .Y(n82) );
  BUFX2 U39 ( .A(n62), .Y(n42) );
  INVX1 U40 ( .A(n42), .Y(n81) );
  BUFX2 U41 ( .A(n63), .Y(n43) );
  INVX1 U42 ( .A(n43), .Y(n80) );
  BUFX2 U43 ( .A(n64), .Y(n44) );
  INVX1 U44 ( .A(n44), .Y(n79) );
  BUFX2 U45 ( .A(n65), .Y(n45) );
  INVX1 U46 ( .A(n45), .Y(n78) );
  BUFX2 U47 ( .A(n66), .Y(n46) );
  INVX1 U48 ( .A(n46), .Y(n77) );
  BUFX2 U49 ( .A(n67), .Y(n47) );
  INVX1 U50 ( .A(n47), .Y(n76) );
  BUFX2 U51 ( .A(n68), .Y(n48) );
  INVX1 U52 ( .A(n48), .Y(n75) );
endmodule


module reg16_20 ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n1, n18, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82;

  dff_362 d0 ( .q(\read<0> ), .d(n82), .clk(clk), .rst(rst) );
  dff_361 d1 ( .q(\read<1> ), .d(n81), .clk(clk), .rst(rst) );
  dff_360 d2 ( .q(\read<2> ), .d(n80), .clk(clk), .rst(rst) );
  dff_359 d3 ( .q(\read<3> ), .d(n79), .clk(clk), .rst(rst) );
  dff_358 d4 ( .q(\read<4> ), .d(n78), .clk(clk), .rst(rst) );
  dff_357 d5 ( .q(\read<5> ), .d(n77), .clk(clk), .rst(rst) );
  dff_356 d6 ( .q(\read<6> ), .d(n76), .clk(clk), .rst(rst) );
  dff_355 d7 ( .q(\read<7> ), .d(n75), .clk(clk), .rst(rst) );
  dff_354 d8 ( .q(\read<8> ), .d(n74), .clk(clk), .rst(rst) );
  dff_353 d9 ( .q(\read<9> ), .d(n73), .clk(clk), .rst(rst) );
  dff_352 d10 ( .q(\read<10> ), .d(n72), .clk(clk), .rst(rst) );
  dff_351 d11 ( .q(\read<11> ), .d(n71), .clk(clk), .rst(rst) );
  dff_350 d12 ( .q(\read<12> ), .d(n70), .clk(clk), .rst(rst) );
  dff_349 d13 ( .q(\read<13> ), .d(n69), .clk(clk), .rst(rst) );
  dff_348 d14 ( .q(\read<14> ), .d(n68), .clk(clk), .rst(rst) );
  dff_347 d15 ( .q(\read<15> ), .d(n67), .clk(clk), .rst(rst) );
  AOI22X1 U18 ( .A(\read<9> ), .B(n49), .C(\write<9> ), .D(wr_en), .Y(n66) );
  AOI22X1 U19 ( .A(\read<8> ), .B(n49), .C(\write<8> ), .D(wr_en), .Y(n65) );
  AOI22X1 U20 ( .A(\read<7> ), .B(n49), .C(\write<7> ), .D(wr_en), .Y(n64) );
  AOI22X1 U21 ( .A(\read<6> ), .B(n49), .C(\write<6> ), .D(wr_en), .Y(n63) );
  AOI22X1 U22 ( .A(\read<5> ), .B(n50), .C(\write<5> ), .D(wr_en), .Y(n62) );
  AOI22X1 U23 ( .A(\read<4> ), .B(n50), .C(\write<4> ), .D(wr_en), .Y(n61) );
  AOI22X1 U24 ( .A(\read<3> ), .B(n50), .C(\write<3> ), .D(wr_en), .Y(n60) );
  AOI22X1 U25 ( .A(\read<2> ), .B(n50), .C(\write<2> ), .D(wr_en), .Y(n59) );
  AOI22X1 U26 ( .A(\read<1> ), .B(n50), .C(\write<1> ), .D(wr_en), .Y(n58) );
  AOI22X1 U27 ( .A(\read<15> ), .B(n50), .C(\write<15> ), .D(wr_en), .Y(n57)
         );
  AOI22X1 U28 ( .A(\read<14> ), .B(n50), .C(\write<14> ), .D(wr_en), .Y(n56)
         );
  AOI22X1 U29 ( .A(\read<13> ), .B(n50), .C(\write<13> ), .D(wr_en), .Y(n55)
         );
  AOI22X1 U30 ( .A(\read<12> ), .B(n50), .C(\write<12> ), .D(wr_en), .Y(n54)
         );
  AOI22X1 U31 ( .A(\read<11> ), .B(n50), .C(\write<11> ), .D(wr_en), .Y(n53)
         );
  AOI22X1 U32 ( .A(\read<10> ), .B(n50), .C(\write<10> ), .D(wr_en), .Y(n52)
         );
  AOI22X1 U33 ( .A(\read<0> ), .B(n50), .C(\write<0> ), .D(wr_en), .Y(n51) );
  INVX1 U1 ( .A(wr_en), .Y(n49) );
  INVX1 U2 ( .A(wr_en), .Y(n50) );
  BUFX2 U3 ( .A(n51), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n82) );
  BUFX2 U5 ( .A(n52), .Y(n18) );
  INVX1 U6 ( .A(n18), .Y(n72) );
  BUFX2 U7 ( .A(n53), .Y(n35) );
  INVX1 U8 ( .A(n35), .Y(n71) );
  BUFX2 U9 ( .A(n54), .Y(n36) );
  INVX1 U10 ( .A(n36), .Y(n70) );
  BUFX2 U11 ( .A(n55), .Y(n37) );
  INVX1 U12 ( .A(n37), .Y(n69) );
  BUFX2 U13 ( .A(n56), .Y(n38) );
  INVX1 U14 ( .A(n38), .Y(n68) );
  BUFX2 U15 ( .A(n57), .Y(n39) );
  INVX1 U16 ( .A(n39), .Y(n67) );
  BUFX2 U17 ( .A(n58), .Y(n40) );
  INVX1 U34 ( .A(n40), .Y(n81) );
  BUFX2 U35 ( .A(n59), .Y(n41) );
  INVX1 U36 ( .A(n41), .Y(n80) );
  BUFX2 U37 ( .A(n60), .Y(n42) );
  INVX1 U38 ( .A(n42), .Y(n79) );
  BUFX2 U39 ( .A(n61), .Y(n43) );
  INVX1 U40 ( .A(n43), .Y(n78) );
  BUFX2 U41 ( .A(n62), .Y(n44) );
  INVX1 U42 ( .A(n44), .Y(n77) );
  BUFX2 U43 ( .A(n63), .Y(n45) );
  INVX1 U44 ( .A(n45), .Y(n76) );
  BUFX2 U45 ( .A(n64), .Y(n46) );
  INVX1 U46 ( .A(n46), .Y(n75) );
  BUFX2 U47 ( .A(n65), .Y(n47) );
  INVX1 U48 ( .A(n47), .Y(n74) );
  BUFX2 U49 ( .A(n66), .Y(n48) );
  INVX1 U50 ( .A(n48), .Y(n73) );
endmodule


module reg16_19 ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n1, n18, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84;

  dff_346 d0 ( .q(\read<0> ), .d(n84), .clk(clk), .rst(rst) );
  dff_345 d1 ( .q(\read<1> ), .d(n83), .clk(clk), .rst(rst) );
  dff_344 d2 ( .q(\read<2> ), .d(n82), .clk(clk), .rst(rst) );
  dff_343 d3 ( .q(\read<3> ), .d(n81), .clk(clk), .rst(rst) );
  dff_342 d4 ( .q(\read<4> ), .d(n80), .clk(clk), .rst(rst) );
  dff_341 d5 ( .q(\read<5> ), .d(n79), .clk(clk), .rst(rst) );
  dff_340 d6 ( .q(\read<6> ), .d(n78), .clk(clk), .rst(rst) );
  dff_339 d7 ( .q(\read<7> ), .d(n77), .clk(clk), .rst(rst) );
  dff_338 d8 ( .q(\read<8> ), .d(n76), .clk(clk), .rst(rst) );
  dff_337 d9 ( .q(\read<9> ), .d(n75), .clk(clk), .rst(rst) );
  dff_336 d10 ( .q(\read<10> ), .d(n74), .clk(clk), .rst(rst) );
  dff_335 d11 ( .q(\read<11> ), .d(n73), .clk(clk), .rst(rst) );
  dff_334 d12 ( .q(\read<12> ), .d(n72), .clk(clk), .rst(rst) );
  dff_333 d13 ( .q(\read<13> ), .d(n71), .clk(clk), .rst(rst) );
  dff_332 d14 ( .q(\read<14> ), .d(n70), .clk(clk), .rst(rst) );
  dff_331 d15 ( .q(\read<15> ), .d(n69), .clk(clk), .rst(rst) );
  AOI22X1 U18 ( .A(\read<9> ), .B(n49), .C(\write<9> ), .D(n50), .Y(n68) );
  AOI22X1 U19 ( .A(\read<8> ), .B(n49), .C(\write<8> ), .D(n50), .Y(n67) );
  AOI22X1 U20 ( .A(\read<7> ), .B(n49), .C(\write<7> ), .D(n50), .Y(n66) );
  AOI22X1 U21 ( .A(\read<6> ), .B(n49), .C(\write<6> ), .D(n50), .Y(n65) );
  AOI22X1 U22 ( .A(\read<5> ), .B(n52), .C(\write<5> ), .D(n50), .Y(n64) );
  AOI22X1 U23 ( .A(\read<4> ), .B(n52), .C(\write<4> ), .D(n50), .Y(n63) );
  AOI22X1 U24 ( .A(\read<3> ), .B(n52), .C(\write<3> ), .D(n50), .Y(n62) );
  AOI22X1 U25 ( .A(\read<2> ), .B(n52), .C(\write<2> ), .D(n50), .Y(n61) );
  AOI22X1 U26 ( .A(\read<1> ), .B(n52), .C(\write<1> ), .D(n50), .Y(n60) );
  AOI22X1 U27 ( .A(\read<15> ), .B(n52), .C(\write<15> ), .D(n50), .Y(n59) );
  AOI22X1 U28 ( .A(\read<14> ), .B(n52), .C(\write<14> ), .D(n50), .Y(n58) );
  AOI22X1 U29 ( .A(\read<13> ), .B(n52), .C(\write<13> ), .D(n50), .Y(n57) );
  AOI22X1 U30 ( .A(\read<12> ), .B(n52), .C(\write<12> ), .D(n51), .Y(n56) );
  AOI22X1 U31 ( .A(\read<11> ), .B(n52), .C(\write<11> ), .D(n51), .Y(n55) );
  AOI22X1 U32 ( .A(\read<10> ), .B(n52), .C(\write<10> ), .D(n51), .Y(n54) );
  AOI22X1 U33 ( .A(\read<0> ), .B(n52), .C(\write<0> ), .D(n51), .Y(n53) );
  INVX1 U1 ( .A(wr_en), .Y(n49) );
  INVX1 U2 ( .A(wr_en), .Y(n52) );
  INVX1 U3 ( .A(n49), .Y(n51) );
  INVX1 U4 ( .A(n49), .Y(n50) );
  BUFX2 U5 ( .A(n53), .Y(n1) );
  INVX1 U6 ( .A(n1), .Y(n84) );
  BUFX2 U7 ( .A(n54), .Y(n18) );
  INVX1 U8 ( .A(n18), .Y(n74) );
  BUFX2 U9 ( .A(n55), .Y(n35) );
  INVX1 U10 ( .A(n35), .Y(n73) );
  BUFX2 U11 ( .A(n56), .Y(n36) );
  INVX1 U12 ( .A(n36), .Y(n72) );
  BUFX2 U13 ( .A(n57), .Y(n37) );
  INVX1 U14 ( .A(n37), .Y(n71) );
  BUFX2 U15 ( .A(n58), .Y(n38) );
  INVX1 U16 ( .A(n38), .Y(n70) );
  BUFX2 U17 ( .A(n59), .Y(n39) );
  INVX1 U34 ( .A(n39), .Y(n69) );
  BUFX2 U35 ( .A(n60), .Y(n40) );
  INVX1 U36 ( .A(n40), .Y(n83) );
  BUFX2 U37 ( .A(n61), .Y(n41) );
  INVX1 U38 ( .A(n41), .Y(n82) );
  BUFX2 U39 ( .A(n62), .Y(n42) );
  INVX1 U40 ( .A(n42), .Y(n81) );
  BUFX2 U41 ( .A(n63), .Y(n43) );
  INVX1 U42 ( .A(n43), .Y(n80) );
  BUFX2 U43 ( .A(n64), .Y(n44) );
  INVX1 U44 ( .A(n44), .Y(n79) );
  BUFX2 U45 ( .A(n65), .Y(n45) );
  INVX1 U46 ( .A(n45), .Y(n78) );
  BUFX2 U47 ( .A(n66), .Y(n46) );
  INVX1 U48 ( .A(n46), .Y(n77) );
  BUFX2 U49 ( .A(n67), .Y(n47) );
  INVX1 U50 ( .A(n47), .Y(n76) );
  BUFX2 U51 ( .A(n68), .Y(n48) );
  INVX1 U52 ( .A(n48), .Y(n75) );
endmodule


module reg1_14 ( d, q, clk, rst, en );
  input d, clk, rst, en;
  output q;
  wire   n1, n2, n3, n4;

  dff_330 d0 ( .q(q), .d(n4), .clk(clk), .rst(rst) );
  INVX1 U1 ( .A(en), .Y(n1) );
  INVX1 U2 ( .A(q), .Y(n3) );
  MUX2X1 U3 ( .B(n2), .A(n3), .S(n1), .Y(n4) );
  INVX1 U4 ( .A(d), .Y(n2) );
endmodule


module reg1_13 ( d, q, clk, rst, en );
  input d, clk, rst, en;
  output q;
  wire   n1, n2, n3;

  dff_329 d0 ( .q(q), .d(n3), .clk(clk), .rst(rst) );
  INVX1 U1 ( .A(q), .Y(n2) );
  INVX1 U2 ( .A(d), .Y(n1) );
  MUX2X1 U3 ( .B(n2), .A(n1), .S(en), .Y(n3) );
endmodule


module reg1_12 ( d, q, clk, rst, en );
  input d, clk, rst, en;
  output q;
  wire   n1, n2, n3, n4;

  dff_328 d0 ( .q(q), .d(n4), .clk(clk), .rst(rst) );
  INVX1 U1 ( .A(en), .Y(n1) );
  INVX1 U2 ( .A(q), .Y(n3) );
  MUX2X1 U3 ( .B(n2), .A(n3), .S(n1), .Y(n4) );
  INVX1 U4 ( .A(d), .Y(n2) );
endmodule


module reg1_11 ( d, q, clk, rst, en );
  input d, clk, rst, en;
  output q;
  wire   n1, n2, n3, n4;

  dff_327 d0 ( .q(q), .d(n4), .clk(clk), .rst(rst) );
  INVX1 U1 ( .A(en), .Y(n1) );
  INVX1 U2 ( .A(q), .Y(n3) );
  INVX1 U3 ( .A(d), .Y(n2) );
  MUX2X1 U4 ( .B(n2), .A(n3), .S(n1), .Y(n4) );
endmodule


module reg1_10 ( d, q, clk, rst, en );
  input d, clk, rst, en;
  output q;
  wire   n1, n2, n3, n4, n5, n6, n7;

  dff_326 d0 ( .q(q), .d(n7), .clk(clk), .rst(rst) );
  OR2X1 U1 ( .A(en), .B(n3), .Y(n5) );
  INVX1 U2 ( .A(q), .Y(n3) );
  INVX1 U3 ( .A(n5), .Y(n4) );
  OR2X1 U4 ( .A(n4), .B(en), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
  INVX1 U6 ( .A(d), .Y(n6) );
  AOI21X1 U7 ( .A(n6), .B(n5), .C(n2), .Y(n7) );
endmodule


module reg1_9 ( d, q, clk, rst, en );
  input d, clk, rst, en;
  output q;
  wire   n1, n3, n5, n6;

  dff_325 d0 ( .q(q), .d(n6), .clk(clk), .rst(rst) );
  AOI22X1 U3 ( .A(en), .B(d), .C(q), .D(n3), .Y(n5) );
  INVX1 U1 ( .A(en), .Y(n3) );
  BUFX2 U2 ( .A(n5), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n6) );
endmodule


module reg1_8 ( d, q, clk, rst, en );
  input d, clk, rst, en;
  output q;
  wire   n1, n3, n5, n6;

  dff_324 d0 ( .q(q), .d(n6), .clk(clk), .rst(rst) );
  AOI22X1 U3 ( .A(en), .B(d), .C(q), .D(n3), .Y(n5) );
  INVX1 U1 ( .A(en), .Y(n3) );
  BUFX2 U2 ( .A(n5), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n6) );
endmodule


module reg1_7 ( d, q, clk, rst, en );
  input d, clk, rst, en;
  output q;
  wire   n1, n3, n5, n6;

  dff_323 d0 ( .q(q), .d(n6), .clk(clk), .rst(rst) );
  AOI22X1 U3 ( .A(en), .B(d), .C(q), .D(n3), .Y(n5) );
  INVX1 U1 ( .A(en), .Y(n3) );
  BUFX2 U2 ( .A(n5), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n6) );
endmodule


module reg16_18 ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n1, n18, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84;

  dff_322 d0 ( .q(\read<0> ), .d(n84), .clk(clk), .rst(rst) );
  dff_321 d1 ( .q(\read<1> ), .d(n83), .clk(clk), .rst(rst) );
  dff_320 d2 ( .q(\read<2> ), .d(n82), .clk(clk), .rst(rst) );
  dff_319 d3 ( .q(\read<3> ), .d(n81), .clk(clk), .rst(rst) );
  dff_318 d4 ( .q(\read<4> ), .d(n80), .clk(clk), .rst(rst) );
  dff_317 d5 ( .q(\read<5> ), .d(n79), .clk(clk), .rst(rst) );
  dff_316 d6 ( .q(\read<6> ), .d(n78), .clk(clk), .rst(rst) );
  dff_315 d7 ( .q(\read<7> ), .d(n77), .clk(clk), .rst(rst) );
  dff_314 d8 ( .q(\read<8> ), .d(n76), .clk(clk), .rst(rst) );
  dff_313 d9 ( .q(\read<9> ), .d(n75), .clk(clk), .rst(rst) );
  dff_312 d10 ( .q(\read<10> ), .d(n74), .clk(clk), .rst(rst) );
  dff_311 d11 ( .q(\read<11> ), .d(n73), .clk(clk), .rst(rst) );
  dff_310 d12 ( .q(\read<12> ), .d(n72), .clk(clk), .rst(rst) );
  dff_309 d13 ( .q(\read<13> ), .d(n71), .clk(clk), .rst(rst) );
  dff_308 d14 ( .q(\read<14> ), .d(n70), .clk(clk), .rst(rst) );
  dff_307 d15 ( .q(\read<15> ), .d(n69), .clk(clk), .rst(rst) );
  AOI22X1 U18 ( .A(\read<9> ), .B(n49), .C(\write<9> ), .D(n50), .Y(n68) );
  AOI22X1 U19 ( .A(\read<8> ), .B(n49), .C(\write<8> ), .D(n50), .Y(n67) );
  AOI22X1 U20 ( .A(\read<7> ), .B(n49), .C(\write<7> ), .D(n50), .Y(n66) );
  AOI22X1 U21 ( .A(\read<6> ), .B(n49), .C(\write<6> ), .D(n50), .Y(n65) );
  AOI22X1 U22 ( .A(\read<5> ), .B(n52), .C(\write<5> ), .D(n50), .Y(n64) );
  AOI22X1 U23 ( .A(\read<4> ), .B(n52), .C(\write<4> ), .D(n50), .Y(n63) );
  AOI22X1 U24 ( .A(\read<3> ), .B(n52), .C(\write<3> ), .D(n50), .Y(n62) );
  AOI22X1 U25 ( .A(\read<2> ), .B(n52), .C(\write<2> ), .D(n50), .Y(n61) );
  AOI22X1 U26 ( .A(\read<1> ), .B(n52), .C(\write<1> ), .D(n50), .Y(n60) );
  AOI22X1 U27 ( .A(\read<15> ), .B(n52), .C(\write<15> ), .D(n50), .Y(n59) );
  AOI22X1 U28 ( .A(\read<14> ), .B(n52), .C(\write<14> ), .D(n50), .Y(n58) );
  AOI22X1 U29 ( .A(\read<13> ), .B(n52), .C(\write<13> ), .D(n50), .Y(n57) );
  AOI22X1 U30 ( .A(\read<12> ), .B(n52), .C(\write<12> ), .D(n51), .Y(n56) );
  AOI22X1 U31 ( .A(\read<11> ), .B(n52), .C(\write<11> ), .D(n51), .Y(n55) );
  AOI22X1 U32 ( .A(\read<10> ), .B(n52), .C(\write<10> ), .D(n51), .Y(n54) );
  AOI22X1 U33 ( .A(\read<0> ), .B(n52), .C(\write<0> ), .D(n51), .Y(n53) );
  INVX1 U1 ( .A(wr_en), .Y(n49) );
  INVX1 U2 ( .A(wr_en), .Y(n52) );
  INVX1 U3 ( .A(n49), .Y(n51) );
  INVX1 U4 ( .A(n49), .Y(n50) );
  BUFX2 U5 ( .A(n53), .Y(n1) );
  INVX1 U6 ( .A(n1), .Y(n84) );
  BUFX2 U7 ( .A(n54), .Y(n18) );
  INVX1 U8 ( .A(n18), .Y(n74) );
  BUFX2 U9 ( .A(n55), .Y(n35) );
  INVX1 U10 ( .A(n35), .Y(n73) );
  BUFX2 U11 ( .A(n56), .Y(n36) );
  INVX1 U12 ( .A(n36), .Y(n72) );
  BUFX2 U13 ( .A(n57), .Y(n37) );
  INVX1 U14 ( .A(n37), .Y(n71) );
  BUFX2 U15 ( .A(n58), .Y(n38) );
  INVX1 U16 ( .A(n38), .Y(n70) );
  BUFX2 U17 ( .A(n59), .Y(n39) );
  INVX1 U34 ( .A(n39), .Y(n69) );
  BUFX2 U35 ( .A(n60), .Y(n40) );
  INVX1 U36 ( .A(n40), .Y(n83) );
  BUFX2 U37 ( .A(n61), .Y(n41) );
  INVX1 U38 ( .A(n41), .Y(n82) );
  BUFX2 U39 ( .A(n62), .Y(n42) );
  INVX1 U40 ( .A(n42), .Y(n81) );
  BUFX2 U41 ( .A(n63), .Y(n43) );
  INVX1 U42 ( .A(n43), .Y(n80) );
  BUFX2 U43 ( .A(n64), .Y(n44) );
  INVX1 U44 ( .A(n44), .Y(n79) );
  BUFX2 U45 ( .A(n65), .Y(n45) );
  INVX1 U46 ( .A(n45), .Y(n78) );
  BUFX2 U47 ( .A(n66), .Y(n46) );
  INVX1 U48 ( .A(n46), .Y(n77) );
  BUFX2 U49 ( .A(n67), .Y(n47) );
  INVX1 U50 ( .A(n47), .Y(n76) );
  BUFX2 U51 ( .A(n68), .Y(n48) );
  INVX1 U52 ( .A(n48), .Y(n75) );
endmodule


module MEM_control ( MemRead, MemWrite, .opcode({\opcode<4> , \opcode<3> , 
        \opcode<2> , \opcode<1> , \opcode<0> }) );
  input \opcode<4> , \opcode<3> , \opcode<2> , \opcode<1> , \opcode<0> ;
  output MemRead, MemWrite;
  wire   n1, n3, n2, n4, n5, n6;

  NOR3X1 U2 ( .A(n1), .B(\opcode<1> ), .C(n6), .Y(MemRead) );
  NOR2X1 U3 ( .A(n6), .B(n3), .Y(MemWrite) );
  XOR2X1 U4 ( .A(\opcode<1> ), .B(\opcode<0> ), .Y(n3) );
  OR2X1 U1 ( .A(\opcode<3> ), .B(\opcode<2> ), .Y(n2) );
  INVX1 U5 ( .A(n2), .Y(n4) );
  AND2X2 U6 ( .A(n4), .B(\opcode<4> ), .Y(n5) );
  INVX1 U7 ( .A(n5), .Y(n6) );
  INVX1 U8 ( .A(\opcode<0> ), .Y(n1) );
endmodule


module WB_control_1 ( MemtoReg, RegWrite, ld_imm, compareS, btr, writeR7, 
        RegDst, .opcode({\opcode<4> , \opcode<3> , \opcode<2> , \opcode<1> , 
        \opcode<0> }) );
  input \opcode<4> , \opcode<3> , \opcode<2> , \opcode<1> , \opcode<0> ;
  output MemtoReg, RegWrite, ld_imm, compareS, btr, writeR7, RegDst;
  wire   n1, n3, n5, n6, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40;

  BUFX2 U1 ( .A(\opcode<2> ), .Y(n1) );
  AND2X2 U2 ( .A(n3), .B(\opcode<4> ), .Y(ld_imm) );
  INVX1 U3 ( .A(n35), .Y(n3) );
  AND2X2 U4 ( .A(n5), .B(\opcode<4> ), .Y(MemtoReg) );
  INVX1 U5 ( .A(n39), .Y(n5) );
  INVX1 U6 ( .A(\opcode<4> ), .Y(n40) );
  OR2X2 U7 ( .A(n9), .B(n40), .Y(n6) );
  INVX1 U8 ( .A(n6), .Y(compareS) );
  AND2X2 U9 ( .A(\opcode<3> ), .B(\opcode<2> ), .Y(n8) );
  INVX1 U10 ( .A(n8), .Y(n9) );
  OR2X2 U11 ( .A(\opcode<2> ), .B(\opcode<1> ), .Y(n10) );
  INVX1 U12 ( .A(n10), .Y(n11) );
  INVX1 U13 ( .A(n10), .Y(n12) );
  INVX1 U14 ( .A(n10), .Y(n13) );
  AND2X1 U15 ( .A(n29), .B(n28), .Y(n14) );
  INVX1 U16 ( .A(n14), .Y(n15) );
  BUFX2 U17 ( .A(n37), .Y(n16) );
  AND2X2 U18 ( .A(\opcode<0> ), .B(\opcode<3> ), .Y(n17) );
  INVX1 U19 ( .A(n17), .Y(n18) );
  BUFX2 U20 ( .A(n33), .Y(n19) );
  OR2X1 U21 ( .A(n32), .B(n31), .Y(n20) );
  INVX1 U22 ( .A(n20), .Y(n21) );
  AND2X1 U23 ( .A(n28), .B(n27), .Y(n22) );
  INVX1 U24 ( .A(n22), .Y(n23) );
  AND2X1 U25 ( .A(n26), .B(n30), .Y(n24) );
  INVX1 U26 ( .A(n24), .Y(n25) );
  INVX1 U27 ( .A(n38), .Y(n26) );
  BUFX2 U28 ( .A(\opcode<1> ), .Y(n27) );
  BUFX2 U29 ( .A(\opcode<4> ), .Y(n28) );
  INVX1 U30 ( .A(\opcode<3> ), .Y(n38) );
  INVX1 U31 ( .A(n36), .Y(n29) );
  INVX1 U32 ( .A(n1), .Y(n30) );
  INVX1 U33 ( .A(n13), .Y(n34) );
  INVX1 U34 ( .A(\opcode<0> ), .Y(n36) );
  MUX2X1 U35 ( .B(n25), .A(n30), .S(n28), .Y(n32) );
  NAND3X1 U36 ( .A(n27), .B(n1), .C(n38), .Y(n33) );
  OAI21X1 U37 ( .A(n15), .B(n27), .C(n19), .Y(n31) );
  OAI21X1 U38 ( .A(n23), .B(n25), .C(n21), .Y(RegDst) );
  NOR2X1 U39 ( .A(n19), .B(n28), .Y(writeR7) );
  NOR3X1 U40 ( .A(n40), .B(n18), .C(n34), .Y(btr) );
  NAND3X1 U41 ( .A(n36), .B(\opcode<3> ), .C(n12), .Y(n35) );
  NAND3X1 U42 ( .A(n36), .B(n26), .C(n28), .Y(n37) );
  NAND3X1 U43 ( .A(n23), .B(n21), .C(n16), .Y(RegWrite) );
  NAND3X1 U44 ( .A(\opcode<0> ), .B(n38), .C(n11), .Y(n39) );
endmodule


module mf_data ( .rd({\rd<2> , \rd<1> , \rd<0> }), .rs({\rs<2> , \rs<1> , 
        \rs<0> }), regdst, memtoreg, slbi, compareS, btr_cntl, .aluOut({
        \aluOut<15> , \aluOut<14> , \aluOut<13> , \aluOut<12> , \aluOut<11> , 
        \aluOut<10> , \aluOut<9> , \aluOut<8> , \aluOut<7> , \aluOut<6> , 
        \aluOut<5> , \aluOut<4> , \aluOut<3> , \aluOut<2> , \aluOut<1> , 
        \aluOut<0> }), .mem_out({\mem_out<15> , \mem_out<14> , \mem_out<13> , 
        \mem_out<12> , \mem_out<11> , \mem_out<10> , \mem_out<9> , 
        \mem_out<8> , \mem_out<7> , \mem_out<6> , \mem_out<5> , \mem_out<4> , 
        \mem_out<3> , \mem_out<2> , \mem_out<1> , \mem_out<0> }), .alu_out({
        \alu_out<15> , \alu_out<14> , \alu_out<13> , \alu_out<12> , 
        \alu_out<11> , \alu_out<10> , \alu_out<9> , \alu_out<8> , \alu_out<7> , 
        \alu_out<6> , \alu_out<5> , \alu_out<4> , \alu_out<3> , \alu_out<2> , 
        \alu_out<1> , \alu_out<0> }), .imm({\imm<15> , \imm<14> , \imm<13> , 
        \imm<12> , \imm<11> , \imm<10> , \imm<9> , \imm<8> , \imm<7> , 
        \imm<6> , \imm<5> , \imm<4> , \imm<3> , \imm<2> , \imm<1> , \imm<0> }), 
    .writereg({\writereg<2> , \writereg<1> , \writereg<0> }), ofl, zero, N, P, 
        cout, .inst({\inst<15> , \inst<14> , \inst<13> , \inst<12> , 
        \inst<11> , \inst<10> , \inst<9> , \inst<8> , \inst<7> , \inst<6> , 
        \inst<5> , \inst<4> , \inst<3> , \inst<2> , \inst<1> , \inst<0> }), 
        ld_imm, .regwritedata({\regwritedata<15> , \regwritedata<14> , 
        \regwritedata<13> , \regwritedata<12> , \regwritedata<11> , 
        \regwritedata<10> , \regwritedata<9> , \regwritedata<8> , 
        \regwritedata<7> , \regwritedata<6> , \regwritedata<5> , 
        \regwritedata<4> , \regwritedata<3> , \regwritedata<2> , 
        \regwritedata<1> , \regwritedata<0> }) );
  input \rd<2> , \rd<1> , \rd<0> , \rs<2> , \rs<1> , \rs<0> , regdst, memtoreg,
         slbi, compareS, btr_cntl, \aluOut<15> , \aluOut<14> , \aluOut<13> ,
         \aluOut<12> , \aluOut<11> , \aluOut<10> , \aluOut<9> , \aluOut<8> ,
         \aluOut<7> , \aluOut<6> , \aluOut<5> , \aluOut<4> , \aluOut<3> ,
         \aluOut<2> , \aluOut<1> , \aluOut<0> , \mem_out<15> , \mem_out<14> ,
         \mem_out<13> , \mem_out<12> , \mem_out<11> , \mem_out<10> ,
         \mem_out<9> , \mem_out<8> , \mem_out<7> , \mem_out<6> , \mem_out<5> ,
         \mem_out<4> , \mem_out<3> , \mem_out<2> , \mem_out<1> , \mem_out<0> ,
         \alu_out<15> , \alu_out<14> , \alu_out<13> , \alu_out<12> ,
         \alu_out<11> , \alu_out<10> , \alu_out<9> , \alu_out<8> ,
         \alu_out<7> , \alu_out<6> , \alu_out<5> , \alu_out<4> , \alu_out<3> ,
         \alu_out<2> , \alu_out<1> , \alu_out<0> , \imm<15> , \imm<14> ,
         \imm<13> , \imm<12> , \imm<11> , \imm<10> , \imm<9> , \imm<8> ,
         \imm<7> , \imm<6> , \imm<5> , \imm<4> , \imm<3> , \imm<2> , \imm<1> ,
         \imm<0> , ofl, zero, N, P, cout, \inst<15> , \inst<14> , \inst<13> ,
         \inst<12> , \inst<11> , \inst<10> , \inst<9> , \inst<8> , \inst<7> ,
         \inst<6> , \inst<5> , \inst<4> , \inst<3> , \inst<2> , \inst<1> ,
         \inst<0> , ld_imm;
  output \writereg<2> , \writereg<1> , \writereg<0> , \regwritedata<15> ,
         \regwritedata<14> , \regwritedata<13> , \regwritedata<12> ,
         \regwritedata<11> , \regwritedata<10> , \regwritedata<9> ,
         \regwritedata<8> , \regwritedata<7> , \regwritedata<6> ,
         \regwritedata<5> , \regwritedata<4> , \regwritedata<3> ,
         \regwritedata<2> , \regwritedata<1> , \regwritedata<0> ;
  wire   n269, n270, n271, n272, n273, n274, n5, n15, n16, n17, n1, n2, n3, n4,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n35, n37, n39, n41,
         n42, n43, n45, n46, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n131, n132, n133,
         n135, n136, n137, n138, n139, n140, n141, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n188, n189, n191, n193,
         n194, n195, n196, n197, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268;

  AOI22X1 U19 ( .A(regdst), .B(\rd<2> ), .C(\rs<2> ), .D(n5), .Y(n15) );
  AOI22X1 U20 ( .A(\rd<1> ), .B(regdst), .C(\rs<1> ), .D(n5), .Y(n16) );
  AOI22X1 U21 ( .A(\rd<0> ), .B(regdst), .C(\rs<0> ), .D(n5), .Y(n17) );
  INVX4 U2 ( .A(n243), .Y(n259) );
  INVX1 U3 ( .A(\imm<0> ), .Y(n209) );
  INVX1 U4 ( .A(\aluOut<2> ), .Y(n226) );
  INVX1 U5 ( .A(\aluOut<15> ), .Y(n206) );
  INVX1 U6 ( .A(\aluOut<13> ), .Y(n227) );
  INVX1 U7 ( .A(\imm<2> ), .Y(n224) );
  INVX1 U8 ( .A(\aluOut<11> ), .Y(n236) );
  INVX1 U9 ( .A(\mem_out<4> ), .Y(n237) );
  INVX1 U10 ( .A(\mem_out<5> ), .Y(n32) );
  INVX1 U11 ( .A(\aluOut<6> ), .Y(n246) );
  INVX1 U12 ( .A(n206), .Y(n201) );
  INVX1 U13 ( .A(\aluOut<7> ), .Y(n29) );
  INVX4 U14 ( .A(slbi), .Y(n257) );
  INVX1 U15 ( .A(n30), .Y(n1) );
  INVX1 U16 ( .A(n241), .Y(n2) );
  INVX1 U17 ( .A(n2), .Y(n3) );
  INVX1 U18 ( .A(n208), .Y(n4) );
  INVX1 U22 ( .A(n4), .Y(n6) );
  INVX1 U23 ( .A(n156), .Y(n7) );
  INVX1 U24 ( .A(ld_imm), .Y(n8) );
  INVX1 U25 ( .A(n8), .Y(n9) );
  AND2X2 U26 ( .A(n98), .B(n19), .Y(n10) );
  OR2X2 U27 ( .A(n85), .B(n21), .Y(n11) );
  INVX1 U28 ( .A(n11), .Y(n250) );
  INVX2 U29 ( .A(btr_cntl), .Y(n21) );
  INVX2 U30 ( .A(ld_imm), .Y(n19) );
  OAI21X1 U31 ( .A(n13), .B(slbi), .C(n104), .Y(n12) );
  INVX1 U32 ( .A(n12), .Y(n258) );
  INVX4 U33 ( .A(n24), .Y(n136) );
  INVX1 U34 ( .A(n8), .Y(n199) );
  INVX1 U35 ( .A(n18), .Y(n13) );
  INVX1 U36 ( .A(n21), .Y(n14) );
  INVX1 U37 ( .A(n21), .Y(n18) );
  OR2X2 U38 ( .A(memtoreg), .B(slbi), .Y(n106) );
  INVX1 U39 ( .A(memtoreg), .Y(n241) );
  INVX1 U40 ( .A(n195), .Y(n20) );
  INVX1 U41 ( .A(n25), .Y(n200) );
  INVX1 U42 ( .A(n33), .Y(n202) );
  INVX1 U43 ( .A(n22), .Y(n242) );
  NOR3X1 U44 ( .A(n23), .B(n153), .C(n193), .Y(n22) );
  INVX8 U45 ( .A(\aluOut<5> ), .Y(n23) );
  OR2X2 U46 ( .A(n3), .B(n9), .Y(n24) );
  INVX1 U47 ( .A(memtoreg), .Y(n25) );
  INVX1 U48 ( .A(n140), .Y(n27) );
  INVX1 U49 ( .A(n259), .Y(n28) );
  NOR3X1 U50 ( .A(n27), .B(n28), .C(n29), .Y(n26) );
  INVX1 U51 ( .A(n26), .Y(n253) );
  INVX4 U52 ( .A(n33), .Y(n204) );
  BUFX2 U53 ( .A(memtoreg), .Y(n30) );
  OAI21X1 U54 ( .A(n53), .B(n32), .C(n103), .Y(n31) );
  INVX1 U55 ( .A(n31), .Y(n245) );
  AND2X2 U56 ( .A(btr_cntl), .B(n257), .Y(n153) );
  INVX1 U57 ( .A(n243), .Y(n261) );
  AND2X2 U58 ( .A(n14), .B(n259), .Y(n239) );
  OR2X2 U59 ( .A(n11), .B(n243), .Y(n33) );
  OR2X2 U60 ( .A(n30), .B(n246), .Y(n247) );
  OR2X2 U61 ( .A(n51), .B(n35), .Y(\regwritedata<0> ) );
  OR2X2 U62 ( .A(n128), .B(n182), .Y(n35) );
  OR2X2 U63 ( .A(n78), .B(n37), .Y(\regwritedata<14> ) );
  OR2X2 U64 ( .A(n79), .B(n131), .Y(n37) );
  OR2X2 U65 ( .A(n81), .B(n39), .Y(\regwritedata<15> ) );
  OR2X2 U66 ( .A(n132), .B(n80), .Y(n39) );
  OR2X2 U67 ( .A(n62), .B(n41), .Y(\regwritedata<4> ) );
  OR2X2 U68 ( .A(n133), .B(n63), .Y(n41) );
  AND2X2 U69 ( .A(n66), .B(n253), .Y(n42) );
  AND2X2 U70 ( .A(n92), .B(n45), .Y(n43) );
  INVX1 U71 ( .A(n43), .Y(\regwritedata<9> ) );
  AND2X2 U72 ( .A(n93), .B(n91), .Y(n45) );
  AND2X2 U73 ( .A(n158), .B(n48), .Y(n46) );
  INVX1 U74 ( .A(n46), .Y(\regwritedata<12> ) );
  AND2X2 U75 ( .A(n97), .B(n76), .Y(n48) );
  AND2X2 U76 ( .A(n95), .B(n89), .Y(n49) );
  INVX1 U77 ( .A(n49), .Y(n50) );
  AND2X2 U78 ( .A(n201), .B(n135), .Y(n51) );
  AND2X2 U79 ( .A(n154), .B(n20), .Y(n52) );
  OR2X2 U80 ( .A(n9), .B(n25), .Y(n53) );
  INVX1 U81 ( .A(n53), .Y(n54) );
  OR2X2 U82 ( .A(n199), .B(n227), .Y(n55) );
  INVX1 U83 ( .A(n55), .Y(n56) );
  OR2X2 U84 ( .A(n100), .B(n199), .Y(n57) );
  INVX1 U85 ( .A(n57), .Y(n58) );
  AND2X2 U86 ( .A(n19), .B(n188), .Y(n59) );
  AND2X2 U87 ( .A(\imm<3> ), .B(n199), .Y(n60) );
  INVX1 U88 ( .A(n60), .Y(n61) );
  AND2X2 U89 ( .A(\imm<4> ), .B(n207), .Y(n62) );
  AND2X2 U90 ( .A(n203), .B(\aluOut<4> ), .Y(n63) );
  OR2X2 U91 ( .A(n24), .B(n237), .Y(n64) );
  AND2X2 U92 ( .A(\mem_out<7> ), .B(n136), .Y(n65) );
  INVX1 U93 ( .A(n65), .Y(n66) );
  AND2X2 U94 ( .A(\aluOut<7> ), .B(n204), .Y(n67) );
  INVX1 U95 ( .A(n67), .Y(n68) );
  AND2X2 U96 ( .A(\aluOut<5> ), .B(n204), .Y(n69) );
  INVX1 U97 ( .A(n69), .Y(n70) );
  AND2X2 U98 ( .A(\imm<10> ), .B(n207), .Y(n71) );
  INVX1 U99 ( .A(n71), .Y(n72) );
  AND2X2 U100 ( .A(\aluOut<4> ), .B(n202), .Y(n73) );
  INVX1 U101 ( .A(n73), .Y(n74) );
  AND2X2 U102 ( .A(\aluOut<12> ), .B(n203), .Y(n75) );
  INVX1 U103 ( .A(n75), .Y(n76) );
  AND2X2 U104 ( .A(\aluOut<13> ), .B(n205), .Y(n77) );
  AND2X2 U105 ( .A(\aluOut<1> ), .B(n204), .Y(n78) );
  AND2X2 U106 ( .A(\aluOut<14> ), .B(n203), .Y(n79) );
  AND2X2 U107 ( .A(\aluOut<0> ), .B(n135), .Y(n80) );
  AND2X2 U108 ( .A(\aluOut<15> ), .B(n205), .Y(n81) );
  BUFX2 U109 ( .A(n252), .Y(n82) );
  OR2X2 U110 ( .A(n208), .B(n162), .Y(n83) );
  INVX1 U111 ( .A(n83), .Y(n84) );
  OR2X2 U112 ( .A(compareS), .B(slbi), .Y(n85) );
  INVX1 U113 ( .A(n85), .Y(n86) );
  BUFX2 U114 ( .A(n234), .Y(n87) );
  AND2X2 U115 ( .A(\imm<1> ), .B(ld_imm), .Y(n88) );
  INVX1 U116 ( .A(n88), .Y(n89) );
  AND2X2 U117 ( .A(\aluOut<6> ), .B(n202), .Y(n90) );
  INVX1 U118 ( .A(n90), .Y(n91) );
  BUFX2 U119 ( .A(n255), .Y(n92) );
  BUFX2 U120 ( .A(n256), .Y(n93) );
  AND2X2 U121 ( .A(n155), .B(n241), .Y(n94) );
  INVX1 U122 ( .A(n94), .Y(n95) );
  AND2X2 U123 ( .A(\aluOut<3> ), .B(n204), .Y(n96) );
  INVX1 U124 ( .A(n96), .Y(n97) );
  AND2X2 U125 ( .A(\aluOut<1> ), .B(n196), .Y(n98) );
  AND2X2 U126 ( .A(\mem_out<2> ), .B(n200), .Y(n99) );
  INVX1 U127 ( .A(n99), .Y(n100) );
  AND2X2 U128 ( .A(n18), .B(n86), .Y(n101) );
  INVX1 U129 ( .A(n101), .Y(n102) );
  OR2X2 U130 ( .A(n243), .B(n242), .Y(n103) );
  AND2X2 U131 ( .A(\aluOut<10> ), .B(n188), .Y(n104) );
  BUFX2 U132 ( .A(n223), .Y(n105) );
  INVX1 U133 ( .A(n106), .Y(n107) );
  AND2X2 U134 ( .A(n160), .B(n24), .Y(n108) );
  INVX1 U135 ( .A(n108), .Y(n109) );
  AND2X2 U136 ( .A(\aluOut<8> ), .B(n205), .Y(n110) );
  INVX1 U137 ( .A(n110), .Y(n111) );
  AND2X2 U138 ( .A(\aluOut<2> ), .B(n204), .Y(n112) );
  INVX1 U139 ( .A(n112), .Y(n113) );
  OR2X2 U140 ( .A(n102), .B(n200), .Y(n114) );
  INVX1 U141 ( .A(n114), .Y(n115) );
  BUFX2 U142 ( .A(n216), .Y(n116) );
  BUFX2 U143 ( .A(n222), .Y(n117) );
  AND2X2 U144 ( .A(\imm<5> ), .B(n251), .Y(n118) );
  INVX1 U145 ( .A(n118), .Y(n119) );
  AND2X2 U146 ( .A(\imm<6> ), .B(n251), .Y(n120) );
  INVX1 U147 ( .A(n120), .Y(n121) );
  OR2X2 U148 ( .A(n247), .B(n7), .Y(n122) );
  INVX1 U149 ( .A(n122), .Y(n123) );
  BUFX2 U150 ( .A(n248), .Y(n124) );
  BUFX2 U151 ( .A(n229), .Y(n125) );
  AND2X2 U152 ( .A(n261), .B(n221), .Y(n126) );
  INVX1 U153 ( .A(n126), .Y(n127) );
  INVX1 U154 ( .A(n219), .Y(n128) );
  AND2X2 U155 ( .A(n82), .B(n42), .Y(n129) );
  INVX1 U156 ( .A(n129), .Y(\regwritedata<7> ) );
  INVX1 U157 ( .A(n266), .Y(n131) );
  INVX1 U158 ( .A(n268), .Y(n132) );
  INVX1 U159 ( .A(n240), .Y(n133) );
  BUFX2 U160 ( .A(compareS), .Y(n208) );
  BUFX2 U161 ( .A(n269), .Y(\regwritedata<13> ) );
  AND2X2 U162 ( .A(n250), .B(n261), .Y(n135) );
  INVX1 U163 ( .A(n260), .Y(n137) );
  INVX1 U164 ( .A(n137), .Y(n138) );
  BUFX2 U165 ( .A(n263), .Y(n139) );
  AND2X2 U166 ( .A(n20), .B(n156), .Y(n140) );
  INVX1 U167 ( .A(n274), .Y(n141) );
  INVX1 U168 ( .A(n141), .Y(\regwritedata<5> ) );
  INVX1 U169 ( .A(n215), .Y(n143) );
  INVX1 U170 ( .A(n143), .Y(n144) );
  OR2X2 U171 ( .A(n200), .B(n209), .Y(n145) );
  INVX1 U172 ( .A(n145), .Y(n146) );
  OR2X2 U173 ( .A(n153), .B(n226), .Y(n147) );
  INVX1 U174 ( .A(n147), .Y(n148) );
  INVX1 U175 ( .A(n254), .Y(n149) );
  INVX1 U176 ( .A(n149), .Y(n150) );
  INVX1 U177 ( .A(n262), .Y(n151) );
  INVX1 U178 ( .A(n151), .Y(n152) );
  INVX1 U179 ( .A(regdst), .Y(n5) );
  INVX1 U180 ( .A(n153), .Y(n154) );
  AND2X1 U181 ( .A(\imm<1> ), .B(slbi), .Y(n155) );
  INVX1 U182 ( .A(n153), .Y(n156) );
  INVX1 U183 ( .A(n264), .Y(n157) );
  INVX1 U184 ( .A(n157), .Y(n158) );
  INVX1 U185 ( .A(n225), .Y(n159) );
  INVX1 U186 ( .A(n159), .Y(n160) );
  AND2X2 U187 ( .A(\aluOut<14> ), .B(n257), .Y(n161) );
  INVX1 U188 ( .A(n161), .Y(n162) );
  INVX1 U189 ( .A(n232), .Y(n163) );
  INVX1 U190 ( .A(n163), .Y(n164) );
  INVX1 U191 ( .A(n64), .Y(n165) );
  INVX1 U192 ( .A(n249), .Y(n166) );
  INVX1 U193 ( .A(n166), .Y(n167) );
  BUFX2 U194 ( .A(n17), .Y(n168) );
  INVX1 U195 ( .A(n168), .Y(\writereg<0> ) );
  BUFX2 U196 ( .A(n16), .Y(n169) );
  INVX1 U197 ( .A(n169), .Y(\writereg<1> ) );
  BUFX2 U198 ( .A(n15), .Y(n170) );
  INVX1 U199 ( .A(n170), .Y(\writereg<2> ) );
  BUFX2 U200 ( .A(n217), .Y(n171) );
  INVX1 U201 ( .A(n235), .Y(n172) );
  INVX1 U202 ( .A(n172), .Y(n173) );
  BUFX2 U203 ( .A(n212), .Y(n174) );
  INVX1 U204 ( .A(n228), .Y(n175) );
  INVX1 U205 ( .A(n175), .Y(n176) );
  INVX1 U206 ( .A(n231), .Y(n177) );
  INVX1 U207 ( .A(n177), .Y(n178) );
  INVX1 U208 ( .A(n77), .Y(n179) );
  INVX1 U209 ( .A(n265), .Y(n180) );
  INVX1 U210 ( .A(n180), .Y(n181) );
  INVX1 U211 ( .A(n220), .Y(n182) );
  INVX1 U212 ( .A(n230), .Y(n183) );
  INVX1 U213 ( .A(n183), .Y(n184) );
  BUFX2 U214 ( .A(n244), .Y(n185) );
  INVX1 U215 ( .A(n272), .Y(n186) );
  INVX1 U216 ( .A(n186), .Y(\regwritedata<8> ) );
  INVX1 U217 ( .A(n195), .Y(n188) );
  INVX1 U218 ( .A(n270), .Y(n189) );
  INVX1 U219 ( .A(n189), .Y(\regwritedata<11> ) );
  INVX1 U220 ( .A(n271), .Y(n191) );
  INVX1 U221 ( .A(n191), .Y(\regwritedata<10> ) );
  INVX1 U222 ( .A(n194), .Y(n193) );
  INVX1 U223 ( .A(n195), .Y(n194) );
  AND2X2 U224 ( .A(compareS), .B(n257), .Y(n195) );
  INVX1 U225 ( .A(n195), .Y(n196) );
  INVX1 U226 ( .A(n273), .Y(n197) );
  INVX1 U227 ( .A(n197), .Y(\regwritedata<6> ) );
  AND2X2 U228 ( .A(n261), .B(n52), .Y(n203) );
  AND2X2 U229 ( .A(n259), .B(n52), .Y(n205) );
  BUFX4 U230 ( .A(n267), .Y(n207) );
  OR2X2 U231 ( .A(memtoreg), .B(ld_imm), .Y(n243) );
  NAND3X1 U232 ( .A(n52), .B(n259), .C(\aluOut<0> ), .Y(n220) );
  AND2X2 U233 ( .A(\inst<15> ), .B(\inst<14> ), .Y(n210) );
  NAND3X1 U234 ( .A(n6), .B(\inst<13> ), .C(n210), .Y(n217) );
  AOI21X1 U235 ( .A(P), .B(\inst<12> ), .C(zero), .Y(n212) );
  MUX2X1 U236 ( .B(P), .A(cout), .S(\inst<12> ), .Y(n211) );
  MUX2X1 U237 ( .B(n174), .A(n211), .S(\inst<11> ), .Y(n213) );
  NAND3X1 U238 ( .A(n8), .B(n213), .C(n107), .Y(n216) );
  AND2X2 U239 ( .A(\mem_out<0> ), .B(n2), .Y(n214) );
  AOI22X1 U240 ( .A(\imm<0> ), .B(n199), .C(n19), .D(n214), .Y(n215) );
  OAI21X1 U241 ( .A(n171), .B(n116), .C(n144), .Y(n218) );
  AOI21X1 U242 ( .A(slbi), .B(n146), .C(n218), .Y(n219) );
  NAND3X1 U243 ( .A(n1), .B(n154), .C(n10), .Y(n223) );
  AOI21X1 U244 ( .A(n54), .B(\mem_out<1> ), .C(n50), .Y(n222) );
  AND2X2 U245 ( .A(n18), .B(n84), .Y(n221) );
  NAND3X1 U246 ( .A(n117), .B(n127), .C(n105), .Y(\regwritedata<1> ) );
  AOI21X1 U247 ( .A(n257), .B(n19), .C(n224), .Y(n225) );
  NAND3X1 U248 ( .A(n259), .B(n148), .C(n188), .Y(n229) );
  AOI21X1 U249 ( .A(n56), .B(n115), .C(n58), .Y(n228) );
  NAND3X1 U250 ( .A(n109), .B(n125), .C(n176), .Y(\regwritedata<2> ) );
  NAND3X1 U251 ( .A(n59), .B(n1), .C(\aluOut<3> ), .Y(n235) );
  AND2X2 U252 ( .A(n86), .B(\aluOut<12> ), .Y(n233) );
  NAND3X1 U253 ( .A(\imm<3> ), .B(n3), .C(slbi), .Y(n231) );
  NAND3X1 U254 ( .A(n19), .B(\mem_out<3> ), .C(n200), .Y(n230) );
  NAND3X1 U255 ( .A(n61), .B(n178), .C(n184), .Y(n232) );
  AOI21X1 U256 ( .A(n239), .B(n233), .C(n164), .Y(n234) );
  OAI21X1 U257 ( .A(n173), .B(n7), .C(n87), .Y(\regwritedata<3> ) );
  OAI21X1 U258 ( .A(n257), .B(n30), .C(n19), .Y(n267) );
  NOR3X1 U259 ( .A(slbi), .B(n6), .C(n236), .Y(n238) );
  AOI21X1 U260 ( .A(n239), .B(n238), .C(n165), .Y(n240) );
  OAI21X1 U261 ( .A(n257), .B(n30), .C(n19), .Y(n251) );
  NAND3X1 U262 ( .A(n250), .B(\aluOut<10> ), .C(n259), .Y(n244) );
  NAND3X1 U263 ( .A(n245), .B(n119), .C(n185), .Y(n274) );
  NAND3X1 U264 ( .A(n259), .B(n250), .C(\aluOut<9> ), .Y(n249) );
  AOI22X1 U265 ( .A(\mem_out<6> ), .B(n136), .C(n59), .D(n123), .Y(n248) );
  NAND3X1 U266 ( .A(n167), .B(n121), .C(n124), .Y(n273) );
  AOI22X1 U267 ( .A(\imm<7> ), .B(n251), .C(\aluOut<8> ), .D(n204), .Y(n252)
         );
  AOI22X1 U268 ( .A(\imm<8> ), .B(n207), .C(\mem_out<8> ), .D(n136), .Y(n254)
         );
  NAND3X1 U269 ( .A(n111), .B(n68), .C(n150), .Y(n272) );
  NAND3X1 U270 ( .A(n140), .B(n259), .C(\aluOut<9> ), .Y(n256) );
  AOI22X1 U271 ( .A(\imm<9> ), .B(n207), .C(\mem_out<9> ), .D(n136), .Y(n255)
         );
  AOI22X1 U272 ( .A(n259), .B(n258), .C(\mem_out<10> ), .D(n136), .Y(n260) );
  NAND3X1 U273 ( .A(n138), .B(n70), .C(n72), .Y(n271) );
  NAND3X1 U274 ( .A(n140), .B(n259), .C(\aluOut<11> ), .Y(n263) );
  AOI22X1 U275 ( .A(\imm<11> ), .B(n251), .C(\mem_out<11> ), .D(n136), .Y(n262) );
  NAND3X1 U276 ( .A(n139), .B(n152), .C(n74), .Y(n270) );
  AOI22X1 U277 ( .A(\imm<12> ), .B(n207), .C(\mem_out<12> ), .D(n136), .Y(n264) );
  AOI22X1 U278 ( .A(\imm<13> ), .B(n207), .C(\mem_out<13> ), .D(n136), .Y(n265) );
  NAND3X1 U279 ( .A(n113), .B(n179), .C(n181), .Y(n269) );
  AOI22X1 U280 ( .A(\imm<14> ), .B(n207), .C(\mem_out<14> ), .D(n136), .Y(n266) );
  AOI22X1 U281 ( .A(\imm<15> ), .B(n207), .C(\mem_out<15> ), .D(n136), .Y(n268) );
endmodule


module reg3_2 ( .read({\read<2> , \read<1> , \read<0> }), .write({\write<2> , 
        \write<1> , \write<0> }), wr_en, rst, clk );
  input \write<2> , \write<1> , \write<0> , wr_en, rst, clk;
  output \read<2> , \read<1> , \read<0> ;
  wire   n1, n5, n9, n10, n11, n12, n13, n14, n15, n16;

  dff_306 d0 ( .q(\read<0> ), .d(n16), .clk(clk), .rst(rst) );
  dff_305 d1 ( .q(\read<1> ), .d(n15), .clk(clk), .rst(rst) );
  dff_304 d2 ( .q(\read<2> ), .d(n14), .clk(clk), .rst(rst) );
  AOI22X1 U5 ( .A(\read<2> ), .B(n10), .C(\write<2> ), .D(wr_en), .Y(n13) );
  AOI22X1 U6 ( .A(\read<1> ), .B(n10), .C(\write<1> ), .D(wr_en), .Y(n12) );
  AOI22X1 U7 ( .A(\read<0> ), .B(n10), .C(\write<0> ), .D(wr_en), .Y(n11) );
  INVX1 U1 ( .A(wr_en), .Y(n10) );
  BUFX2 U2 ( .A(n11), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(n16) );
  BUFX2 U4 ( .A(n12), .Y(n5) );
  INVX1 U8 ( .A(n5), .Y(n15) );
  BUFX2 U9 ( .A(n13), .Y(n9) );
  INVX1 U10 ( .A(n9), .Y(n14) );
endmodule


module reg3_1 ( .read({\read<2> , \read<1> , \read<0> }), .write({\write<2> , 
        \write<1> , \write<0> }), wr_en, rst, clk );
  input \write<2> , \write<1> , \write<0> , wr_en, rst, clk;
  output \read<2> , \read<1> , \read<0> ;
  wire   n1, n5, n9, n10, n11, n12, n13, n14, n15, n16;

  dff_303 d0 ( .q(\read<0> ), .d(n16), .clk(clk), .rst(rst) );
  dff_302 d1 ( .q(\read<1> ), .d(n15), .clk(clk), .rst(rst) );
  dff_301 d2 ( .q(\read<2> ), .d(n14), .clk(clk), .rst(rst) );
  AOI22X1 U5 ( .A(\read<2> ), .B(n10), .C(\write<2> ), .D(wr_en), .Y(n13) );
  AOI22X1 U6 ( .A(\read<1> ), .B(n10), .C(\write<1> ), .D(wr_en), .Y(n12) );
  AOI22X1 U7 ( .A(\read<0> ), .B(n10), .C(\write<0> ), .D(wr_en), .Y(n11) );
  INVX1 U1 ( .A(wr_en), .Y(n10) );
  BUFX2 U2 ( .A(n11), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(n16) );
  BUFX2 U4 ( .A(n12), .Y(n5) );
  INVX1 U8 ( .A(n5), .Y(n15) );
  BUFX2 U9 ( .A(n13), .Y(n9) );
  INVX1 U10 ( .A(n9), .Y(n14) );
endmodule


module reg3_0 ( .read({\read<2> , \read<1> , \read<0> }), .write({\write<2> , 
        \write<1> , \write<0> }), wr_en, rst, clk );
  input \write<2> , \write<1> , \write<0> , wr_en, rst, clk;
  output \read<2> , \read<1> , \read<0> ;
  wire   n1, n5, n9, n10, n11, n12, n13, n14, n15, n16;

  dff_300 d0 ( .q(\read<0> ), .d(n16), .clk(clk), .rst(rst) );
  dff_299 d1 ( .q(\read<1> ), .d(n15), .clk(clk), .rst(rst) );
  dff_298 d2 ( .q(\read<2> ), .d(n14), .clk(clk), .rst(rst) );
  AOI22X1 U5 ( .A(\read<2> ), .B(n10), .C(\write<2> ), .D(wr_en), .Y(n13) );
  AOI22X1 U6 ( .A(\read<1> ), .B(n10), .C(\write<1> ), .D(wr_en), .Y(n12) );
  AOI22X1 U7 ( .A(\read<0> ), .B(n10), .C(\write<0> ), .D(wr_en), .Y(n11) );
  INVX1 U1 ( .A(wr_en), .Y(n10) );
  BUFX2 U2 ( .A(n11), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(n16) );
  BUFX2 U4 ( .A(n12), .Y(n5) );
  INVX1 U8 ( .A(n5), .Y(n15) );
  BUFX2 U9 ( .A(n13), .Y(n9) );
  INVX1 U10 ( .A(n9), .Y(n14) );
endmodule


module reg16_17 ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n1, n18, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89;

  dff_297 d0 ( .q(\read<0> ), .d(n89), .clk(clk), .rst(rst) );
  dff_296 d1 ( .q(\read<1> ), .d(n88), .clk(clk), .rst(rst) );
  dff_295 d2 ( .q(\read<2> ), .d(n87), .clk(clk), .rst(rst) );
  dff_294 d3 ( .q(\read<3> ), .d(n86), .clk(clk), .rst(rst) );
  dff_293 d4 ( .q(\read<4> ), .d(n85), .clk(clk), .rst(rst) );
  dff_292 d5 ( .q(\read<5> ), .d(n84), .clk(clk), .rst(rst) );
  dff_291 d6 ( .q(\read<6> ), .d(n83), .clk(clk), .rst(rst) );
  dff_290 d7 ( .q(\read<7> ), .d(n82), .clk(clk), .rst(rst) );
  dff_289 d8 ( .q(\read<8> ), .d(n81), .clk(clk), .rst(rst) );
  dff_288 d9 ( .q(\read<9> ), .d(n80), .clk(clk), .rst(rst) );
  dff_287 d10 ( .q(\read<10> ), .d(n79), .clk(clk), .rst(rst) );
  dff_286 d11 ( .q(\read<11> ), .d(n78), .clk(clk), .rst(rst) );
  dff_285 d12 ( .q(\read<12> ), .d(n77), .clk(clk), .rst(rst) );
  dff_284 d13 ( .q(\read<13> ), .d(n76), .clk(clk), .rst(rst) );
  dff_283 d14 ( .q(\read<14> ), .d(n75), .clk(clk), .rst(rst) );
  dff_282 d15 ( .q(\read<15> ), .d(n74), .clk(clk), .rst(rst) );
  AOI22X1 U18 ( .A(\read<9> ), .B(n54), .C(\write<9> ), .D(n55), .Y(n73) );
  AOI22X1 U19 ( .A(\read<8> ), .B(n54), .C(\write<8> ), .D(n55), .Y(n72) );
  AOI22X1 U20 ( .A(\read<7> ), .B(n54), .C(\write<7> ), .D(n55), .Y(n71) );
  AOI22X1 U21 ( .A(\read<6> ), .B(n54), .C(\write<6> ), .D(n55), .Y(n70) );
  AOI22X1 U22 ( .A(\read<5> ), .B(n57), .C(\write<5> ), .D(n55), .Y(n69) );
  AOI22X1 U23 ( .A(\read<4> ), .B(n57), .C(\write<4> ), .D(n55), .Y(n68) );
  AOI22X1 U24 ( .A(\read<3> ), .B(n57), .C(\write<3> ), .D(n55), .Y(n67) );
  AOI22X1 U25 ( .A(\read<2> ), .B(n57), .C(\write<2> ), .D(n55), .Y(n66) );
  AOI22X1 U26 ( .A(\read<1> ), .B(n57), .C(\write<1> ), .D(n55), .Y(n65) );
  AOI22X1 U27 ( .A(n50), .B(n57), .C(\write<15> ), .D(n55), .Y(n64) );
  AOI22X1 U28 ( .A(n53), .B(n57), .C(\write<14> ), .D(n55), .Y(n63) );
  AOI22X1 U29 ( .A(n52), .B(n57), .C(\write<13> ), .D(n55), .Y(n62) );
  AOI22X1 U30 ( .A(n49), .B(n57), .C(\write<12> ), .D(n56), .Y(n61) );
  AOI22X1 U31 ( .A(n51), .B(n57), .C(\write<11> ), .D(n56), .Y(n60) );
  AOI22X1 U32 ( .A(\read<10> ), .B(n57), .C(\write<10> ), .D(n56), .Y(n59) );
  AOI22X1 U33 ( .A(\read<0> ), .B(n57), .C(\write<0> ), .D(n56), .Y(n58) );
  INVX1 U1 ( .A(wr_en), .Y(n54) );
  INVX1 U2 ( .A(wr_en), .Y(n57) );
  INVX1 U3 ( .A(n54), .Y(n56) );
  INVX1 U4 ( .A(n54), .Y(n55) );
  BUFX2 U5 ( .A(n58), .Y(n1) );
  INVX1 U6 ( .A(n1), .Y(n89) );
  BUFX2 U7 ( .A(n59), .Y(n18) );
  INVX1 U8 ( .A(n18), .Y(n79) );
  BUFX2 U9 ( .A(n60), .Y(n35) );
  INVX1 U10 ( .A(n35), .Y(n78) );
  BUFX2 U11 ( .A(n61), .Y(n36) );
  INVX1 U12 ( .A(n36), .Y(n77) );
  BUFX2 U13 ( .A(n62), .Y(n37) );
  INVX1 U14 ( .A(n37), .Y(n76) );
  BUFX2 U15 ( .A(n63), .Y(n38) );
  INVX1 U16 ( .A(n38), .Y(n75) );
  BUFX2 U17 ( .A(n64), .Y(n39) );
  INVX1 U34 ( .A(n39), .Y(n74) );
  BUFX2 U35 ( .A(n65), .Y(n40) );
  INVX1 U36 ( .A(n40), .Y(n88) );
  BUFX2 U37 ( .A(n66), .Y(n41) );
  INVX1 U38 ( .A(n41), .Y(n87) );
  BUFX2 U39 ( .A(n67), .Y(n42) );
  INVX1 U40 ( .A(n42), .Y(n86) );
  BUFX2 U41 ( .A(n68), .Y(n43) );
  INVX1 U42 ( .A(n43), .Y(n85) );
  BUFX2 U43 ( .A(n69), .Y(n44) );
  INVX1 U44 ( .A(n44), .Y(n84) );
  BUFX2 U45 ( .A(n70), .Y(n45) );
  INVX1 U46 ( .A(n45), .Y(n83) );
  BUFX2 U47 ( .A(n71), .Y(n46) );
  INVX1 U48 ( .A(n46), .Y(n82) );
  BUFX2 U49 ( .A(n72), .Y(n47) );
  INVX1 U50 ( .A(n47), .Y(n81) );
  BUFX2 U51 ( .A(n73), .Y(n48) );
  INVX1 U52 ( .A(n48), .Y(n80) );
  BUFX2 U53 ( .A(\read<12> ), .Y(n49) );
  BUFX2 U54 ( .A(\read<15> ), .Y(n50) );
  BUFX2 U55 ( .A(\read<11> ), .Y(n51) );
  BUFX2 U56 ( .A(\read<13> ), .Y(n52) );
  BUFX2 U57 ( .A(\read<14> ), .Y(n53) );
endmodule


module reg16_16 ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n1, n18, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83;

  dff_281 d0 ( .q(\read<0> ), .d(n83), .clk(clk), .rst(rst) );
  dff_280 d1 ( .q(\read<1> ), .d(n82), .clk(clk), .rst(rst) );
  dff_279 d2 ( .q(\read<2> ), .d(n81), .clk(clk), .rst(rst) );
  dff_278 d3 ( .q(\read<3> ), .d(n80), .clk(clk), .rst(rst) );
  dff_277 d4 ( .q(\read<4> ), .d(n79), .clk(clk), .rst(rst) );
  dff_276 d5 ( .q(\read<5> ), .d(n78), .clk(clk), .rst(rst) );
  dff_275 d6 ( .q(\read<6> ), .d(n77), .clk(clk), .rst(rst) );
  dff_274 d7 ( .q(\read<7> ), .d(n76), .clk(clk), .rst(rst) );
  dff_273 d8 ( .q(\read<8> ), .d(n75), .clk(clk), .rst(rst) );
  dff_272 d9 ( .q(\read<9> ), .d(n74), .clk(clk), .rst(rst) );
  dff_271 d10 ( .q(\read<10> ), .d(n73), .clk(clk), .rst(rst) );
  dff_270 d11 ( .q(\read<11> ), .d(n72), .clk(clk), .rst(rst) );
  dff_269 d12 ( .q(\read<12> ), .d(n71), .clk(clk), .rst(rst) );
  dff_268 d13 ( .q(\read<13> ), .d(n70), .clk(clk), .rst(rst) );
  dff_267 d14 ( .q(\read<14> ), .d(n69), .clk(clk), .rst(rst) );
  dff_266 d15 ( .q(\read<15> ), .d(n68), .clk(clk), .rst(rst) );
  AOI22X1 U18 ( .A(\read<9> ), .B(n49), .C(\write<9> ), .D(n50), .Y(n67) );
  AOI22X1 U19 ( .A(\read<8> ), .B(n49), .C(\write<8> ), .D(n50), .Y(n66) );
  AOI22X1 U20 ( .A(\read<7> ), .B(n49), .C(\write<7> ), .D(n50), .Y(n65) );
  AOI22X1 U21 ( .A(\read<6> ), .B(n49), .C(\write<6> ), .D(n50), .Y(n64) );
  AOI22X1 U22 ( .A(\read<5> ), .B(n51), .C(\write<5> ), .D(n50), .Y(n63) );
  AOI22X1 U23 ( .A(\read<4> ), .B(n51), .C(\write<4> ), .D(n50), .Y(n62) );
  AOI22X1 U24 ( .A(\read<3> ), .B(n51), .C(\write<3> ), .D(n50), .Y(n61) );
  AOI22X1 U25 ( .A(\read<2> ), .B(n51), .C(\write<2> ), .D(n50), .Y(n60) );
  AOI22X1 U26 ( .A(\read<1> ), .B(n51), .C(\write<1> ), .D(n50), .Y(n59) );
  AOI22X1 U27 ( .A(\read<15> ), .B(n51), .C(\write<15> ), .D(n50), .Y(n58) );
  AOI22X1 U28 ( .A(\read<14> ), .B(n51), .C(\write<14> ), .D(n50), .Y(n57) );
  AOI22X1 U29 ( .A(\read<13> ), .B(n51), .C(\write<13> ), .D(n50), .Y(n56) );
  AOI22X1 U30 ( .A(\read<12> ), .B(n51), .C(\write<12> ), .D(wr_en), .Y(n55)
         );
  AOI22X1 U31 ( .A(\read<11> ), .B(n51), .C(\write<11> ), .D(wr_en), .Y(n54)
         );
  AOI22X1 U32 ( .A(\read<10> ), .B(n51), .C(\write<10> ), .D(wr_en), .Y(n53)
         );
  AOI22X1 U33 ( .A(\read<0> ), .B(n51), .C(\write<0> ), .D(wr_en), .Y(n52) );
  INVX1 U1 ( .A(wr_en), .Y(n49) );
  INVX1 U2 ( .A(wr_en), .Y(n51) );
  INVX1 U3 ( .A(n49), .Y(n50) );
  BUFX2 U4 ( .A(n52), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n83) );
  BUFX2 U6 ( .A(n53), .Y(n18) );
  INVX1 U7 ( .A(n18), .Y(n73) );
  BUFX2 U8 ( .A(n54), .Y(n35) );
  INVX1 U9 ( .A(n35), .Y(n72) );
  BUFX2 U10 ( .A(n55), .Y(n36) );
  INVX1 U11 ( .A(n36), .Y(n71) );
  BUFX2 U12 ( .A(n56), .Y(n37) );
  INVX1 U13 ( .A(n37), .Y(n70) );
  BUFX2 U14 ( .A(n57), .Y(n38) );
  INVX1 U15 ( .A(n38), .Y(n69) );
  BUFX2 U16 ( .A(n58), .Y(n39) );
  INVX1 U17 ( .A(n39), .Y(n68) );
  BUFX2 U34 ( .A(n59), .Y(n40) );
  INVX1 U35 ( .A(n40), .Y(n82) );
  BUFX2 U36 ( .A(n60), .Y(n41) );
  INVX1 U37 ( .A(n41), .Y(n81) );
  BUFX2 U38 ( .A(n61), .Y(n42) );
  INVX1 U39 ( .A(n42), .Y(n80) );
  BUFX2 U40 ( .A(n62), .Y(n43) );
  INVX1 U41 ( .A(n43), .Y(n79) );
  BUFX2 U42 ( .A(n63), .Y(n44) );
  INVX1 U43 ( .A(n44), .Y(n78) );
  BUFX2 U44 ( .A(n64), .Y(n45) );
  INVX1 U45 ( .A(n45), .Y(n77) );
  BUFX2 U46 ( .A(n65), .Y(n46) );
  INVX1 U47 ( .A(n46), .Y(n76) );
  BUFX2 U48 ( .A(n66), .Y(n47) );
  INVX1 U49 ( .A(n47), .Y(n75) );
  BUFX2 U50 ( .A(n67), .Y(n48) );
  INVX1 U51 ( .A(n48), .Y(n74) );
endmodule


module reg16_15 ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n1, n18, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81;

  dff_265 d0 ( .q(\read<0> ), .d(n81), .clk(clk), .rst(rst) );
  dff_264 d1 ( .q(\read<1> ), .d(n80), .clk(clk), .rst(rst) );
  dff_263 d2 ( .q(\read<2> ), .d(n79), .clk(clk), .rst(rst) );
  dff_262 d3 ( .q(\read<3> ), .d(n78), .clk(clk), .rst(rst) );
  dff_261 d4 ( .q(\read<4> ), .d(n77), .clk(clk), .rst(rst) );
  dff_260 d5 ( .q(\read<5> ), .d(n76), .clk(clk), .rst(rst) );
  dff_259 d6 ( .q(\read<6> ), .d(n75), .clk(clk), .rst(rst) );
  dff_258 d7 ( .q(\read<7> ), .d(n74), .clk(clk), .rst(rst) );
  dff_257 d8 ( .q(\read<8> ), .d(n73), .clk(clk), .rst(rst) );
  dff_256 d9 ( .q(\read<9> ), .d(n72), .clk(clk), .rst(rst) );
  dff_255 d10 ( .q(\read<10> ), .d(n71), .clk(clk), .rst(rst) );
  dff_254 d11 ( .q(\read<11> ), .d(n70), .clk(clk), .rst(rst) );
  dff_253 d12 ( .q(\read<12> ), .d(n69), .clk(clk), .rst(rst) );
  dff_252 d13 ( .q(\read<13> ), .d(n68), .clk(clk), .rst(rst) );
  dff_251 d14 ( .q(\read<14> ), .d(n67), .clk(clk), .rst(rst) );
  dff_250 d15 ( .q(\read<15> ), .d(n66), .clk(clk), .rst(rst) );
  AOI22X1 U18 ( .A(\read<9> ), .B(n49), .C(\write<9> ), .D(wr_en), .Y(n65) );
  AOI22X1 U19 ( .A(\read<8> ), .B(n49), .C(\write<8> ), .D(wr_en), .Y(n64) );
  AOI22X1 U20 ( .A(\read<7> ), .B(n49), .C(\write<7> ), .D(wr_en), .Y(n63) );
  AOI22X1 U21 ( .A(\read<6> ), .B(n49), .C(\write<6> ), .D(wr_en), .Y(n62) );
  AOI22X1 U22 ( .A(\read<5> ), .B(n49), .C(\write<5> ), .D(wr_en), .Y(n61) );
  AOI22X1 U23 ( .A(\read<4> ), .B(n49), .C(\write<4> ), .D(wr_en), .Y(n60) );
  AOI22X1 U24 ( .A(\read<3> ), .B(n49), .C(\write<3> ), .D(wr_en), .Y(n59) );
  AOI22X1 U25 ( .A(\read<2> ), .B(n49), .C(\write<2> ), .D(wr_en), .Y(n58) );
  AOI22X1 U26 ( .A(\read<1> ), .B(n49), .C(\write<1> ), .D(wr_en), .Y(n57) );
  AOI22X1 U27 ( .A(\read<15> ), .B(n49), .C(\write<15> ), .D(wr_en), .Y(n56)
         );
  AOI22X1 U28 ( .A(\read<14> ), .B(n49), .C(\write<14> ), .D(wr_en), .Y(n55)
         );
  AOI22X1 U29 ( .A(\read<13> ), .B(n49), .C(\write<13> ), .D(wr_en), .Y(n54)
         );
  AOI22X1 U30 ( .A(\read<12> ), .B(n49), .C(\write<12> ), .D(wr_en), .Y(n53)
         );
  AOI22X1 U31 ( .A(\read<11> ), .B(n49), .C(\write<11> ), .D(wr_en), .Y(n52)
         );
  AOI22X1 U32 ( .A(\read<10> ), .B(n49), .C(\write<10> ), .D(wr_en), .Y(n51)
         );
  AOI22X1 U33 ( .A(\read<0> ), .B(n49), .C(\write<0> ), .D(wr_en), .Y(n50) );
  INVX1 U1 ( .A(wr_en), .Y(n49) );
  BUFX2 U2 ( .A(n50), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(n81) );
  BUFX2 U4 ( .A(n51), .Y(n18) );
  INVX1 U5 ( .A(n18), .Y(n71) );
  BUFX2 U6 ( .A(n52), .Y(n35) );
  INVX1 U7 ( .A(n35), .Y(n70) );
  BUFX2 U8 ( .A(n53), .Y(n36) );
  INVX1 U9 ( .A(n36), .Y(n69) );
  BUFX2 U10 ( .A(n54), .Y(n37) );
  INVX1 U11 ( .A(n37), .Y(n68) );
  BUFX2 U12 ( .A(n55), .Y(n38) );
  INVX1 U13 ( .A(n38), .Y(n67) );
  BUFX2 U14 ( .A(n56), .Y(n39) );
  INVX1 U15 ( .A(n39), .Y(n66) );
  BUFX2 U16 ( .A(n57), .Y(n40) );
  INVX1 U17 ( .A(n40), .Y(n80) );
  BUFX2 U34 ( .A(n58), .Y(n41) );
  INVX1 U35 ( .A(n41), .Y(n79) );
  BUFX2 U36 ( .A(n59), .Y(n42) );
  INVX1 U37 ( .A(n42), .Y(n78) );
  BUFX2 U38 ( .A(n60), .Y(n43) );
  INVX1 U39 ( .A(n43), .Y(n77) );
  BUFX2 U40 ( .A(n61), .Y(n44) );
  INVX1 U41 ( .A(n44), .Y(n76) );
  BUFX2 U42 ( .A(n62), .Y(n45) );
  INVX1 U43 ( .A(n45), .Y(n75) );
  BUFX2 U44 ( .A(n63), .Y(n46) );
  INVX1 U45 ( .A(n46), .Y(n74) );
  BUFX2 U46 ( .A(n64), .Y(n47) );
  INVX1 U47 ( .A(n47), .Y(n73) );
  BUFX2 U48 ( .A(n65), .Y(n48) );
  INVX1 U49 ( .A(n48), .Y(n72) );
endmodule


module reg16_14 ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n1, n18, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83;

  dff_249 d0 ( .q(\read<0> ), .d(n83), .clk(clk), .rst(rst) );
  dff_248 d1 ( .q(\read<1> ), .d(n82), .clk(clk), .rst(rst) );
  dff_247 d2 ( .q(\read<2> ), .d(n81), .clk(clk), .rst(rst) );
  dff_246 d3 ( .q(\read<3> ), .d(n80), .clk(clk), .rst(rst) );
  dff_245 d4 ( .q(\read<4> ), .d(n79), .clk(clk), .rst(rst) );
  dff_244 d5 ( .q(\read<5> ), .d(n78), .clk(clk), .rst(rst) );
  dff_243 d6 ( .q(\read<6> ), .d(n77), .clk(clk), .rst(rst) );
  dff_242 d7 ( .q(\read<7> ), .d(n76), .clk(clk), .rst(rst) );
  dff_241 d8 ( .q(\read<8> ), .d(n75), .clk(clk), .rst(rst) );
  dff_240 d9 ( .q(\read<9> ), .d(n74), .clk(clk), .rst(rst) );
  dff_239 d10 ( .q(\read<10> ), .d(n73), .clk(clk), .rst(rst) );
  dff_238 d11 ( .q(\read<11> ), .d(n72), .clk(clk), .rst(rst) );
  dff_237 d12 ( .q(\read<12> ), .d(n71), .clk(clk), .rst(rst) );
  dff_236 d13 ( .q(\read<13> ), .d(n70), .clk(clk), .rst(rst) );
  dff_235 d14 ( .q(\read<14> ), .d(n69), .clk(clk), .rst(rst) );
  dff_234 d15 ( .q(\read<15> ), .d(n68), .clk(clk), .rst(rst) );
  AOI22X1 U18 ( .A(\read<9> ), .B(n49), .C(\write<9> ), .D(n50), .Y(n67) );
  AOI22X1 U19 ( .A(\read<8> ), .B(n49), .C(\write<8> ), .D(n50), .Y(n66) );
  AOI22X1 U20 ( .A(\read<7> ), .B(n49), .C(\write<7> ), .D(n50), .Y(n65) );
  AOI22X1 U21 ( .A(\read<6> ), .B(n49), .C(\write<6> ), .D(n50), .Y(n64) );
  AOI22X1 U22 ( .A(\read<5> ), .B(n51), .C(\write<5> ), .D(n50), .Y(n63) );
  AOI22X1 U23 ( .A(\read<4> ), .B(n51), .C(\write<4> ), .D(n50), .Y(n62) );
  AOI22X1 U24 ( .A(\read<3> ), .B(n51), .C(\write<3> ), .D(n50), .Y(n61) );
  AOI22X1 U25 ( .A(\read<2> ), .B(n51), .C(\write<2> ), .D(n50), .Y(n60) );
  AOI22X1 U26 ( .A(\read<1> ), .B(n51), .C(\write<1> ), .D(n50), .Y(n59) );
  AOI22X1 U27 ( .A(\read<15> ), .B(n51), .C(\write<15> ), .D(n50), .Y(n58) );
  AOI22X1 U28 ( .A(\read<14> ), .B(n51), .C(\write<14> ), .D(n50), .Y(n57) );
  AOI22X1 U29 ( .A(\read<13> ), .B(n51), .C(\write<13> ), .D(n50), .Y(n56) );
  AOI22X1 U30 ( .A(\read<12> ), .B(n51), .C(\write<12> ), .D(wr_en), .Y(n55)
         );
  AOI22X1 U31 ( .A(\read<11> ), .B(n51), .C(\write<11> ), .D(wr_en), .Y(n54)
         );
  AOI22X1 U32 ( .A(\read<10> ), .B(n51), .C(\write<10> ), .D(wr_en), .Y(n53)
         );
  AOI22X1 U33 ( .A(\read<0> ), .B(n51), .C(\write<0> ), .D(wr_en), .Y(n52) );
  INVX1 U1 ( .A(wr_en), .Y(n49) );
  INVX1 U2 ( .A(wr_en), .Y(n51) );
  INVX1 U3 ( .A(n49), .Y(n50) );
  BUFX2 U4 ( .A(n52), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n83) );
  BUFX2 U6 ( .A(n53), .Y(n18) );
  INVX1 U7 ( .A(n18), .Y(n73) );
  BUFX2 U8 ( .A(n54), .Y(n35) );
  INVX1 U9 ( .A(n35), .Y(n72) );
  BUFX2 U10 ( .A(n55), .Y(n36) );
  INVX1 U11 ( .A(n36), .Y(n71) );
  BUFX2 U12 ( .A(n56), .Y(n37) );
  INVX1 U13 ( .A(n37), .Y(n70) );
  BUFX2 U14 ( .A(n57), .Y(n38) );
  INVX1 U15 ( .A(n38), .Y(n69) );
  BUFX2 U16 ( .A(n58), .Y(n39) );
  INVX1 U17 ( .A(n39), .Y(n68) );
  BUFX2 U34 ( .A(n59), .Y(n40) );
  INVX1 U35 ( .A(n40), .Y(n82) );
  BUFX2 U36 ( .A(n60), .Y(n41) );
  INVX1 U37 ( .A(n41), .Y(n81) );
  BUFX2 U38 ( .A(n61), .Y(n42) );
  INVX1 U39 ( .A(n42), .Y(n80) );
  BUFX2 U40 ( .A(n62), .Y(n43) );
  INVX1 U41 ( .A(n43), .Y(n79) );
  BUFX2 U42 ( .A(n63), .Y(n44) );
  INVX1 U43 ( .A(n44), .Y(n78) );
  BUFX2 U44 ( .A(n64), .Y(n45) );
  INVX1 U45 ( .A(n45), .Y(n77) );
  BUFX2 U46 ( .A(n65), .Y(n46) );
  INVX1 U47 ( .A(n46), .Y(n76) );
  BUFX2 U48 ( .A(n66), .Y(n47) );
  INVX1 U49 ( .A(n47), .Y(n75) );
  BUFX2 U50 ( .A(n67), .Y(n48) );
  INVX1 U51 ( .A(n48), .Y(n74) );
endmodule


module reg16_13 ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n1, n18, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81;

  dff_233 d0 ( .q(\read<0> ), .d(n81), .clk(clk), .rst(rst) );
  dff_232 d1 ( .q(\read<1> ), .d(n80), .clk(clk), .rst(rst) );
  dff_231 d2 ( .q(\read<2> ), .d(n79), .clk(clk), .rst(rst) );
  dff_230 d3 ( .q(\read<3> ), .d(n78), .clk(clk), .rst(rst) );
  dff_229 d4 ( .q(\read<4> ), .d(n77), .clk(clk), .rst(rst) );
  dff_228 d5 ( .q(\read<5> ), .d(n76), .clk(clk), .rst(rst) );
  dff_227 d6 ( .q(\read<6> ), .d(n75), .clk(clk), .rst(rst) );
  dff_226 d7 ( .q(\read<7> ), .d(n74), .clk(clk), .rst(rst) );
  dff_225 d8 ( .q(\read<8> ), .d(n73), .clk(clk), .rst(rst) );
  dff_224 d9 ( .q(\read<9> ), .d(n72), .clk(clk), .rst(rst) );
  dff_223 d10 ( .q(\read<10> ), .d(n71), .clk(clk), .rst(rst) );
  dff_222 d11 ( .q(\read<11> ), .d(n70), .clk(clk), .rst(rst) );
  dff_221 d12 ( .q(\read<12> ), .d(n69), .clk(clk), .rst(rst) );
  dff_220 d13 ( .q(\read<13> ), .d(n68), .clk(clk), .rst(rst) );
  dff_219 d14 ( .q(\read<14> ), .d(n67), .clk(clk), .rst(rst) );
  dff_218 d15 ( .q(\read<15> ), .d(n66), .clk(clk), .rst(rst) );
  AOI22X1 U18 ( .A(\read<9> ), .B(n49), .C(\write<9> ), .D(wr_en), .Y(n65) );
  AOI22X1 U19 ( .A(\read<8> ), .B(n49), .C(\write<8> ), .D(wr_en), .Y(n64) );
  AOI22X1 U20 ( .A(\read<7> ), .B(n49), .C(\write<7> ), .D(wr_en), .Y(n63) );
  AOI22X1 U21 ( .A(\read<6> ), .B(n49), .C(\write<6> ), .D(wr_en), .Y(n62) );
  AOI22X1 U22 ( .A(\read<5> ), .B(n49), .C(\write<5> ), .D(wr_en), .Y(n61) );
  AOI22X1 U23 ( .A(\read<4> ), .B(n49), .C(\write<4> ), .D(wr_en), .Y(n60) );
  AOI22X1 U24 ( .A(\read<3> ), .B(n49), .C(\write<3> ), .D(wr_en), .Y(n59) );
  AOI22X1 U25 ( .A(\read<2> ), .B(n49), .C(\write<2> ), .D(wr_en), .Y(n58) );
  AOI22X1 U26 ( .A(\read<1> ), .B(n49), .C(\write<1> ), .D(wr_en), .Y(n57) );
  AOI22X1 U27 ( .A(\read<15> ), .B(n49), .C(\write<15> ), .D(wr_en), .Y(n56)
         );
  AOI22X1 U28 ( .A(\read<14> ), .B(n49), .C(\write<14> ), .D(wr_en), .Y(n55)
         );
  AOI22X1 U29 ( .A(\read<13> ), .B(n49), .C(\write<13> ), .D(wr_en), .Y(n54)
         );
  AOI22X1 U30 ( .A(\read<12> ), .B(n49), .C(\write<12> ), .D(wr_en), .Y(n53)
         );
  AOI22X1 U31 ( .A(\read<11> ), .B(n49), .C(\write<11> ), .D(wr_en), .Y(n52)
         );
  AOI22X1 U32 ( .A(\read<10> ), .B(n49), .C(\write<10> ), .D(wr_en), .Y(n51)
         );
  AOI22X1 U33 ( .A(\read<0> ), .B(n49), .C(\write<0> ), .D(wr_en), .Y(n50) );
  INVX1 U1 ( .A(wr_en), .Y(n49) );
  BUFX2 U2 ( .A(n50), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(n81) );
  BUFX2 U4 ( .A(n51), .Y(n18) );
  INVX1 U5 ( .A(n18), .Y(n71) );
  BUFX2 U6 ( .A(n52), .Y(n35) );
  INVX1 U7 ( .A(n35), .Y(n70) );
  BUFX2 U8 ( .A(n53), .Y(n36) );
  INVX1 U9 ( .A(n36), .Y(n69) );
  BUFX2 U10 ( .A(n54), .Y(n37) );
  INVX1 U11 ( .A(n37), .Y(n68) );
  BUFX2 U12 ( .A(n55), .Y(n38) );
  INVX1 U13 ( .A(n38), .Y(n67) );
  BUFX2 U14 ( .A(n56), .Y(n39) );
  INVX1 U15 ( .A(n39), .Y(n66) );
  BUFX2 U16 ( .A(n57), .Y(n40) );
  INVX1 U17 ( .A(n40), .Y(n80) );
  BUFX2 U34 ( .A(n58), .Y(n41) );
  INVX1 U35 ( .A(n41), .Y(n79) );
  BUFX2 U36 ( .A(n59), .Y(n42) );
  INVX1 U37 ( .A(n42), .Y(n78) );
  BUFX2 U38 ( .A(n60), .Y(n43) );
  INVX1 U39 ( .A(n43), .Y(n77) );
  BUFX2 U40 ( .A(n61), .Y(n44) );
  INVX1 U41 ( .A(n44), .Y(n76) );
  BUFX2 U42 ( .A(n62), .Y(n45) );
  INVX1 U43 ( .A(n45), .Y(n75) );
  BUFX2 U44 ( .A(n63), .Y(n46) );
  INVX1 U45 ( .A(n46), .Y(n74) );
  BUFX2 U46 ( .A(n64), .Y(n47) );
  INVX1 U47 ( .A(n47), .Y(n73) );
  BUFX2 U48 ( .A(n65), .Y(n48) );
  INVX1 U49 ( .A(n48), .Y(n72) );
endmodule


module reg16_12 ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n1, n18, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83;

  dff_217 d0 ( .q(\read<0> ), .d(n83), .clk(clk), .rst(rst) );
  dff_216 d1 ( .q(\read<1> ), .d(n82), .clk(clk), .rst(rst) );
  dff_215 d2 ( .q(\read<2> ), .d(n81), .clk(clk), .rst(rst) );
  dff_214 d3 ( .q(\read<3> ), .d(n80), .clk(clk), .rst(rst) );
  dff_213 d4 ( .q(\read<4> ), .d(n79), .clk(clk), .rst(rst) );
  dff_212 d5 ( .q(\read<5> ), .d(n78), .clk(clk), .rst(rst) );
  dff_211 d6 ( .q(\read<6> ), .d(n77), .clk(clk), .rst(rst) );
  dff_210 d7 ( .q(\read<7> ), .d(n76), .clk(clk), .rst(rst) );
  dff_209 d8 ( .q(\read<8> ), .d(n75), .clk(clk), .rst(rst) );
  dff_208 d9 ( .q(\read<9> ), .d(n74), .clk(clk), .rst(rst) );
  dff_207 d10 ( .q(\read<10> ), .d(n73), .clk(clk), .rst(rst) );
  dff_206 d11 ( .q(\read<11> ), .d(n72), .clk(clk), .rst(rst) );
  dff_205 d12 ( .q(\read<12> ), .d(n71), .clk(clk), .rst(rst) );
  dff_204 d13 ( .q(\read<13> ), .d(n70), .clk(clk), .rst(rst) );
  dff_203 d14 ( .q(\read<14> ), .d(n69), .clk(clk), .rst(rst) );
  dff_202 d15 ( .q(\read<15> ), .d(n68), .clk(clk), .rst(rst) );
  AOI22X1 U18 ( .A(\read<9> ), .B(n49), .C(\write<9> ), .D(n50), .Y(n67) );
  AOI22X1 U19 ( .A(\read<8> ), .B(n49), .C(\write<8> ), .D(n50), .Y(n66) );
  AOI22X1 U20 ( .A(\read<7> ), .B(n49), .C(\write<7> ), .D(n50), .Y(n65) );
  AOI22X1 U21 ( .A(\read<6> ), .B(n49), .C(\write<6> ), .D(n50), .Y(n64) );
  AOI22X1 U22 ( .A(\read<5> ), .B(n51), .C(\write<5> ), .D(n50), .Y(n63) );
  AOI22X1 U23 ( .A(\read<4> ), .B(n51), .C(\write<4> ), .D(n50), .Y(n62) );
  AOI22X1 U24 ( .A(\read<3> ), .B(n51), .C(\write<3> ), .D(n50), .Y(n61) );
  AOI22X1 U25 ( .A(\read<2> ), .B(n51), .C(\write<2> ), .D(n50), .Y(n60) );
  AOI22X1 U26 ( .A(\read<1> ), .B(n51), .C(\write<1> ), .D(n50), .Y(n59) );
  AOI22X1 U27 ( .A(\read<15> ), .B(n51), .C(\write<15> ), .D(n50), .Y(n58) );
  AOI22X1 U28 ( .A(\read<14> ), .B(n51), .C(\write<14> ), .D(n50), .Y(n57) );
  AOI22X1 U29 ( .A(\read<13> ), .B(n51), .C(\write<13> ), .D(n50), .Y(n56) );
  AOI22X1 U30 ( .A(\read<12> ), .B(n51), .C(\write<12> ), .D(wr_en), .Y(n55)
         );
  AOI22X1 U31 ( .A(\read<11> ), .B(n51), .C(\write<11> ), .D(wr_en), .Y(n54)
         );
  AOI22X1 U32 ( .A(\read<10> ), .B(n51), .C(\write<10> ), .D(wr_en), .Y(n53)
         );
  AOI22X1 U33 ( .A(\read<0> ), .B(n51), .C(\write<0> ), .D(wr_en), .Y(n52) );
  INVX1 U1 ( .A(wr_en), .Y(n49) );
  INVX1 U2 ( .A(wr_en), .Y(n51) );
  INVX1 U3 ( .A(n49), .Y(n50) );
  BUFX2 U4 ( .A(n52), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n83) );
  BUFX2 U6 ( .A(n53), .Y(n18) );
  INVX1 U7 ( .A(n18), .Y(n73) );
  BUFX2 U8 ( .A(n54), .Y(n35) );
  INVX1 U9 ( .A(n35), .Y(n72) );
  BUFX2 U10 ( .A(n55), .Y(n36) );
  INVX1 U11 ( .A(n36), .Y(n71) );
  BUFX2 U12 ( .A(n56), .Y(n37) );
  INVX1 U13 ( .A(n37), .Y(n70) );
  BUFX2 U14 ( .A(n57), .Y(n38) );
  INVX1 U15 ( .A(n38), .Y(n69) );
  BUFX2 U16 ( .A(n58), .Y(n39) );
  INVX1 U17 ( .A(n39), .Y(n68) );
  BUFX2 U34 ( .A(n59), .Y(n40) );
  INVX1 U35 ( .A(n40), .Y(n82) );
  BUFX2 U36 ( .A(n60), .Y(n41) );
  INVX1 U37 ( .A(n41), .Y(n81) );
  BUFX2 U38 ( .A(n61), .Y(n42) );
  INVX1 U39 ( .A(n42), .Y(n80) );
  BUFX2 U40 ( .A(n62), .Y(n43) );
  INVX1 U41 ( .A(n43), .Y(n79) );
  BUFX2 U42 ( .A(n63), .Y(n44) );
  INVX1 U43 ( .A(n44), .Y(n78) );
  BUFX2 U44 ( .A(n64), .Y(n45) );
  INVX1 U45 ( .A(n45), .Y(n77) );
  BUFX2 U46 ( .A(n65), .Y(n46) );
  INVX1 U47 ( .A(n46), .Y(n76) );
  BUFX2 U48 ( .A(n66), .Y(n47) );
  INVX1 U49 ( .A(n47), .Y(n75) );
  BUFX2 U50 ( .A(n67), .Y(n48) );
  INVX1 U51 ( .A(n48), .Y(n74) );
endmodule


module reg16_11 ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n1, n18, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83;

  dff_201 d0 ( .q(\read<0> ), .d(n83), .clk(clk), .rst(rst) );
  dff_200 d1 ( .q(\read<1> ), .d(n82), .clk(clk), .rst(rst) );
  dff_199 d2 ( .q(\read<2> ), .d(n81), .clk(clk), .rst(rst) );
  dff_198 d3 ( .q(\read<3> ), .d(n80), .clk(clk), .rst(rst) );
  dff_197 d4 ( .q(\read<4> ), .d(n79), .clk(clk), .rst(rst) );
  dff_196 d5 ( .q(\read<5> ), .d(n78), .clk(clk), .rst(rst) );
  dff_195 d6 ( .q(\read<6> ), .d(n77), .clk(clk), .rst(rst) );
  dff_194 d7 ( .q(\read<7> ), .d(n76), .clk(clk), .rst(rst) );
  dff_193 d8 ( .q(\read<8> ), .d(n75), .clk(clk), .rst(rst) );
  dff_192 d9 ( .q(\read<9> ), .d(n74), .clk(clk), .rst(rst) );
  dff_191 d10 ( .q(\read<10> ), .d(n73), .clk(clk), .rst(rst) );
  dff_190 d11 ( .q(\read<11> ), .d(n72), .clk(clk), .rst(rst) );
  dff_189 d12 ( .q(\read<12> ), .d(n71), .clk(clk), .rst(rst) );
  dff_188 d13 ( .q(\read<13> ), .d(n70), .clk(clk), .rst(rst) );
  dff_187 d14 ( .q(\read<14> ), .d(n69), .clk(clk), .rst(rst) );
  dff_186 d15 ( .q(\read<15> ), .d(n68), .clk(clk), .rst(rst) );
  AOI22X1 U18 ( .A(\read<9> ), .B(n49), .C(\write<9> ), .D(n50), .Y(n67) );
  AOI22X1 U19 ( .A(\read<8> ), .B(n49), .C(\write<8> ), .D(n50), .Y(n66) );
  AOI22X1 U20 ( .A(\read<7> ), .B(n49), .C(\write<7> ), .D(n50), .Y(n65) );
  AOI22X1 U21 ( .A(\read<6> ), .B(n49), .C(\write<6> ), .D(n50), .Y(n64) );
  AOI22X1 U22 ( .A(\read<5> ), .B(n51), .C(\write<5> ), .D(n50), .Y(n63) );
  AOI22X1 U23 ( .A(\read<4> ), .B(n51), .C(\write<4> ), .D(n50), .Y(n62) );
  AOI22X1 U24 ( .A(\read<3> ), .B(n51), .C(\write<3> ), .D(n50), .Y(n61) );
  AOI22X1 U25 ( .A(\read<2> ), .B(n51), .C(\write<2> ), .D(n50), .Y(n60) );
  AOI22X1 U26 ( .A(\read<1> ), .B(n51), .C(\write<1> ), .D(n50), .Y(n59) );
  AOI22X1 U27 ( .A(\read<15> ), .B(n51), .C(\write<15> ), .D(n50), .Y(n58) );
  AOI22X1 U28 ( .A(\read<14> ), .B(n51), .C(\write<14> ), .D(n50), .Y(n57) );
  AOI22X1 U29 ( .A(\read<13> ), .B(n51), .C(\write<13> ), .D(n50), .Y(n56) );
  AOI22X1 U30 ( .A(\read<12> ), .B(n51), .C(\write<12> ), .D(wr_en), .Y(n55)
         );
  AOI22X1 U31 ( .A(\read<11> ), .B(n51), .C(\write<11> ), .D(wr_en), .Y(n54)
         );
  AOI22X1 U32 ( .A(\read<10> ), .B(n51), .C(\write<10> ), .D(wr_en), .Y(n53)
         );
  AOI22X1 U33 ( .A(\read<0> ), .B(n51), .C(\write<0> ), .D(wr_en), .Y(n52) );
  INVX1 U1 ( .A(wr_en), .Y(n49) );
  INVX1 U2 ( .A(wr_en), .Y(n51) );
  INVX1 U3 ( .A(n49), .Y(n50) );
  BUFX2 U4 ( .A(n52), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n83) );
  BUFX2 U6 ( .A(n53), .Y(n18) );
  INVX1 U7 ( .A(n18), .Y(n73) );
  BUFX2 U8 ( .A(n54), .Y(n35) );
  INVX1 U9 ( .A(n35), .Y(n72) );
  BUFX2 U10 ( .A(n55), .Y(n36) );
  INVX1 U11 ( .A(n36), .Y(n71) );
  BUFX2 U12 ( .A(n56), .Y(n37) );
  INVX1 U13 ( .A(n37), .Y(n70) );
  BUFX2 U14 ( .A(n57), .Y(n38) );
  INVX1 U15 ( .A(n38), .Y(n69) );
  BUFX2 U16 ( .A(n58), .Y(n39) );
  INVX1 U17 ( .A(n39), .Y(n68) );
  BUFX2 U34 ( .A(n59), .Y(n40) );
  INVX1 U35 ( .A(n40), .Y(n82) );
  BUFX2 U36 ( .A(n60), .Y(n41) );
  INVX1 U37 ( .A(n41), .Y(n81) );
  BUFX2 U38 ( .A(n61), .Y(n42) );
  INVX1 U39 ( .A(n42), .Y(n80) );
  BUFX2 U40 ( .A(n62), .Y(n43) );
  INVX1 U41 ( .A(n43), .Y(n79) );
  BUFX2 U42 ( .A(n63), .Y(n44) );
  INVX1 U43 ( .A(n44), .Y(n78) );
  BUFX2 U44 ( .A(n64), .Y(n45) );
  INVX1 U45 ( .A(n45), .Y(n77) );
  BUFX2 U46 ( .A(n65), .Y(n46) );
  INVX1 U47 ( .A(n46), .Y(n76) );
  BUFX2 U48 ( .A(n66), .Y(n47) );
  INVX1 U49 ( .A(n47), .Y(n75) );
  BUFX2 U50 ( .A(n67), .Y(n48) );
  INVX1 U51 ( .A(n48), .Y(n74) );
endmodule


module reg1_6 ( d, q, clk, rst, en );
  input d, clk, rst, en;
  output q;
  wire   n1, n3, n5, n6;

  dff_185 d0 ( .q(q), .d(n6), .clk(clk), .rst(rst) );
  AOI22X1 U3 ( .A(en), .B(d), .C(q), .D(n3), .Y(n5) );
  INVX1 U1 ( .A(en), .Y(n3) );
  BUFX2 U2 ( .A(n5), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n6) );
endmodule


module reg1_5 ( d, q, clk, rst, en );
  input d, clk, rst, en;
  output q;
  wire   n1, n3, n5, n6;

  dff_184 d0 ( .q(q), .d(n6), .clk(clk), .rst(rst) );
  AOI22X1 U3 ( .A(en), .B(d), .C(q), .D(n3), .Y(n5) );
  INVX1 U1 ( .A(en), .Y(n3) );
  BUFX2 U2 ( .A(n5), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n6) );
endmodule


module reg1_4 ( d, q, clk, rst, en );
  input d, clk, rst, en;
  output q;
  wire   n1, n3, n5, n6;

  dff_183 d0 ( .q(q), .d(n6), .clk(clk), .rst(rst) );
  AOI22X1 U3 ( .A(en), .B(d), .C(q), .D(n3), .Y(n5) );
  INVX1 U1 ( .A(en), .Y(n3) );
  BUFX2 U2 ( .A(n5), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n6) );
endmodule


module reg1_3 ( d, q, clk, rst, en );
  input d, clk, rst, en;
  output q;
  wire   n1, n3, n5, n6;

  dff_182 d0 ( .q(q), .d(n6), .clk(clk), .rst(rst) );
  AOI22X1 U3 ( .A(en), .B(d), .C(q), .D(n3), .Y(n5) );
  INVX1 U1 ( .A(en), .Y(n3) );
  BUFX2 U2 ( .A(n5), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n6) );
endmodule


module reg1_2 ( d, q, clk, rst, en );
  input d, clk, rst, en;
  output q;
  wire   n1, n3, n5, n6;

  dff_181 d0 ( .q(q), .d(n6), .clk(clk), .rst(rst) );
  AOI22X1 U3 ( .A(en), .B(d), .C(q), .D(n3), .Y(n5) );
  INVX1 U1 ( .A(en), .Y(n3) );
  BUFX2 U2 ( .A(n5), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n6) );
endmodule


module reg1_1 ( d, q, clk, rst, en );
  input d, clk, rst, en;
  output q;
  wire   n1, n3, n5, n6;

  dff_180 d0 ( .q(q), .d(n6), .clk(clk), .rst(rst) );
  AOI22X1 U3 ( .A(en), .B(d), .C(q), .D(n3), .Y(n5) );
  INVX1 U1 ( .A(en), .Y(n3) );
  BUFX2 U2 ( .A(n5), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n6) );
endmodule


module reg1_0 ( d, q, clk, rst, en );
  input d, clk, rst, en;
  output q;
  wire   n1, n3, n5, n6;

  dff_179 d0 ( .q(q), .d(n6), .clk(clk), .rst(rst) );
  AOI22X1 U3 ( .A(en), .B(d), .C(q), .D(n3), .Y(n5) );
  INVX1 U1 ( .A(en), .Y(n3) );
  BUFX2 U2 ( .A(n5), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n6) );
endmodule


module reg16_10 ( .read({\read<15> , \read<14> , \read<13> , \read<12> , 
        \read<11> , \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , 
        \read<5> , \read<4> , \read<3> , \read<2> , \read<1> , \read<0> }), 
    .write({\write<15> , \write<14> , \write<13> , \write<12> , \write<11> , 
        \write<10> , \write<9> , \write<8> , \write<7> , \write<6> , 
        \write<5> , \write<4> , \write<3> , \write<2> , \write<1> , \write<0> 
        }), wr_en, rst, clk );
  input \write<15> , \write<14> , \write<13> , \write<12> , \write<11> ,
         \write<10> , \write<9> , \write<8> , \write<7> , \write<6> ,
         \write<5> , \write<4> , \write<3> , \write<2> , \write<1> ,
         \write<0> , wr_en, rst, clk;
  output \read<15> , \read<14> , \read<13> , \read<12> , \read<11> ,
         \read<10> , \read<9> , \read<8> , \read<7> , \read<6> , \read<5> ,
         \read<4> , \read<3> , \read<2> , \read<1> , \read<0> ;
  wire   n1, n18, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81;

  dff_178 d0 ( .q(\read<0> ), .d(n81), .clk(clk), .rst(rst) );
  dff_177 d1 ( .q(\read<1> ), .d(n80), .clk(clk), .rst(rst) );
  dff_176 d2 ( .q(\read<2> ), .d(n79), .clk(clk), .rst(rst) );
  dff_175 d3 ( .q(\read<3> ), .d(n78), .clk(clk), .rst(rst) );
  dff_174 d4 ( .q(\read<4> ), .d(n77), .clk(clk), .rst(rst) );
  dff_173 d5 ( .q(\read<5> ), .d(n76), .clk(clk), .rst(rst) );
  dff_172 d6 ( .q(\read<6> ), .d(n75), .clk(clk), .rst(rst) );
  dff_171 d7 ( .q(\read<7> ), .d(n74), .clk(clk), .rst(rst) );
  dff_170 d8 ( .q(\read<8> ), .d(n73), .clk(clk), .rst(rst) );
  dff_169 d9 ( .q(\read<9> ), .d(n72), .clk(clk), .rst(rst) );
  dff_168 d10 ( .q(\read<10> ), .d(n71), .clk(clk), .rst(rst) );
  dff_167 d11 ( .q(\read<11> ), .d(n70), .clk(clk), .rst(rst) );
  dff_166 d12 ( .q(\read<12> ), .d(n69), .clk(clk), .rst(rst) );
  dff_165 d13 ( .q(\read<13> ), .d(n68), .clk(clk), .rst(rst) );
  dff_164 d14 ( .q(\read<14> ), .d(n67), .clk(clk), .rst(rst) );
  dff_163 d15 ( .q(\read<15> ), .d(n66), .clk(clk), .rst(rst) );
  AOI22X1 U18 ( .A(\read<9> ), .B(n49), .C(\write<9> ), .D(wr_en), .Y(n65) );
  AOI22X1 U19 ( .A(\read<8> ), .B(n49), .C(\write<8> ), .D(wr_en), .Y(n64) );
  AOI22X1 U20 ( .A(\read<7> ), .B(n49), .C(\write<7> ), .D(wr_en), .Y(n63) );
  AOI22X1 U21 ( .A(\read<6> ), .B(n49), .C(\write<6> ), .D(wr_en), .Y(n62) );
  AOI22X1 U22 ( .A(\read<5> ), .B(n49), .C(\write<5> ), .D(wr_en), .Y(n61) );
  AOI22X1 U23 ( .A(\read<4> ), .B(n49), .C(\write<4> ), .D(wr_en), .Y(n60) );
  AOI22X1 U24 ( .A(\read<3> ), .B(n49), .C(\write<3> ), .D(wr_en), .Y(n59) );
  AOI22X1 U25 ( .A(\read<2> ), .B(n49), .C(\write<2> ), .D(wr_en), .Y(n58) );
  AOI22X1 U26 ( .A(\read<1> ), .B(n49), .C(\write<1> ), .D(wr_en), .Y(n57) );
  AOI22X1 U27 ( .A(\read<15> ), .B(n49), .C(\write<15> ), .D(wr_en), .Y(n56)
         );
  AOI22X1 U28 ( .A(\read<14> ), .B(n49), .C(\write<14> ), .D(wr_en), .Y(n55)
         );
  AOI22X1 U29 ( .A(\read<13> ), .B(n49), .C(\write<13> ), .D(wr_en), .Y(n54)
         );
  AOI22X1 U30 ( .A(\read<12> ), .B(n49), .C(\write<12> ), .D(wr_en), .Y(n53)
         );
  AOI22X1 U31 ( .A(\read<11> ), .B(n49), .C(\write<11> ), .D(wr_en), .Y(n52)
         );
  AOI22X1 U32 ( .A(\read<10> ), .B(n49), .C(\write<10> ), .D(wr_en), .Y(n51)
         );
  AOI22X1 U33 ( .A(\read<0> ), .B(n49), .C(\write<0> ), .D(wr_en), .Y(n50) );
  INVX1 U1 ( .A(wr_en), .Y(n49) );
  BUFX2 U2 ( .A(n50), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(n81) );
  BUFX2 U4 ( .A(n51), .Y(n18) );
  INVX1 U5 ( .A(n18), .Y(n71) );
  BUFX2 U6 ( .A(n52), .Y(n35) );
  INVX1 U7 ( .A(n35), .Y(n70) );
  BUFX2 U8 ( .A(n53), .Y(n36) );
  INVX1 U9 ( .A(n36), .Y(n69) );
  BUFX2 U10 ( .A(n54), .Y(n37) );
  INVX1 U11 ( .A(n37), .Y(n68) );
  BUFX2 U12 ( .A(n55), .Y(n38) );
  INVX1 U13 ( .A(n38), .Y(n67) );
  BUFX2 U14 ( .A(n56), .Y(n39) );
  INVX1 U15 ( .A(n39), .Y(n66) );
  BUFX2 U16 ( .A(n57), .Y(n40) );
  INVX1 U17 ( .A(n40), .Y(n80) );
  BUFX2 U34 ( .A(n58), .Y(n41) );
  INVX1 U35 ( .A(n41), .Y(n79) );
  BUFX2 U36 ( .A(n59), .Y(n42) );
  INVX1 U37 ( .A(n42), .Y(n78) );
  BUFX2 U38 ( .A(n60), .Y(n43) );
  INVX1 U39 ( .A(n43), .Y(n77) );
  BUFX2 U40 ( .A(n61), .Y(n44) );
  INVX1 U41 ( .A(n44), .Y(n76) );
  BUFX2 U42 ( .A(n62), .Y(n45) );
  INVX1 U43 ( .A(n45), .Y(n75) );
  BUFX2 U44 ( .A(n63), .Y(n46) );
  INVX1 U45 ( .A(n46), .Y(n74) );
  BUFX2 U46 ( .A(n64), .Y(n47) );
  INVX1 U47 ( .A(n47), .Y(n73) );
  BUFX2 U48 ( .A(n65), .Y(n48) );
  INVX1 U49 ( .A(n48), .Y(n72) );
endmodule


module WB_control_0 ( MemtoReg, RegWrite, ld_imm, compareS, btr, writeR7, 
        RegDst, .opcode({\opcode<4> , \opcode<3> , \opcode<2> , \opcode<1> , 
        \opcode<0> }) );
  input \opcode<4> , \opcode<3> , \opcode<2> , \opcode<1> , \opcode<0> ;
  output MemtoReg, RegWrite, ld_imm, compareS, btr, writeR7, RegDst;
  wire   n1, n2, n3, n4, n5, n6, n8, n9, n10, n11, n12, n14, n16, n18, n19,
         n20, n21, n22, n23, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53;

  INVX2 U1 ( .A(n12), .Y(btr) );
  OR2X1 U2 ( .A(n32), .B(n25), .Y(RegWrite) );
  INVX1 U3 ( .A(n36), .Y(n1) );
  NOR3X1 U4 ( .A(n6), .B(n5), .C(n8), .Y(n2) );
  INVX1 U5 ( .A(\opcode<1> ), .Y(n3) );
  INVX1 U6 ( .A(n3), .Y(n4) );
  INVX4 U7 ( .A(n14), .Y(compareS) );
  INVX1 U8 ( .A(n37), .Y(n5) );
  INVX1 U9 ( .A(\opcode<3> ), .Y(n6) );
  AND2X2 U10 ( .A(n20), .B(n2), .Y(ld_imm) );
  AND2X1 U11 ( .A(n42), .B(n3), .Y(n20) );
  INVX1 U12 ( .A(n51), .Y(n8) );
  INVX1 U13 ( .A(\opcode<3> ), .Y(n9) );
  INVX1 U14 ( .A(n9), .Y(n10) );
  OR2X2 U15 ( .A(\opcode<2> ), .B(\opcode<1> ), .Y(n18) );
  INVX1 U16 ( .A(\opcode<2> ), .Y(n11) );
  AND2X2 U17 ( .A(n51), .B(n50), .Y(n26) );
  OR2X2 U18 ( .A(n21), .B(n18), .Y(n12) );
  OR2X2 U19 ( .A(n23), .B(n49), .Y(n14) );
  OR2X2 U20 ( .A(n19), .B(n38), .Y(n16) );
  INVX1 U21 ( .A(n16), .Y(MemtoReg) );
  BUFX2 U22 ( .A(n53), .Y(n19) );
  BUFX2 U23 ( .A(n48), .Y(n21) );
  AND2X2 U24 ( .A(\opcode<2> ), .B(\opcode<3> ), .Y(n22) );
  INVX1 U25 ( .A(n22), .Y(n23) );
  OR2X1 U26 ( .A(n26), .B(n30), .Y(n25) );
  INVX1 U27 ( .A(n35), .Y(n50) );
  BUFX2 U28 ( .A(n43), .Y(n27) );
  AND2X1 U29 ( .A(n40), .B(n39), .Y(n28) );
  INVX1 U30 ( .A(n28), .Y(n29) );
  OR2X1 U31 ( .A(n45), .B(n44), .Y(n30) );
  INVX1 U32 ( .A(n30), .Y(n31) );
  AND2X1 U33 ( .A(n1), .B(n40), .Y(n32) );
  INVX1 U34 ( .A(n32), .Y(n33) );
  AND2X1 U35 ( .A(n41), .B(n42), .Y(n34) );
  INVX1 U36 ( .A(n34), .Y(n35) );
  AND2X2 U37 ( .A(n6), .B(n36), .Y(n46) );
  INVX1 U38 ( .A(\opcode<4> ), .Y(n36) );
  INVX1 U39 ( .A(n36), .Y(n37) );
  OR2X2 U40 ( .A(n10), .B(\opcode<2> ), .Y(n38) );
  INVX1 U41 ( .A(n11), .Y(n39) );
  INVX1 U42 ( .A(n52), .Y(n40) );
  INVX1 U43 ( .A(n6), .Y(n41) );
  INVX1 U44 ( .A(\opcode<0> ), .Y(n51) );
  INVX1 U45 ( .A(\opcode<2> ), .Y(n42) );
  INVX1 U46 ( .A(\opcode<1> ), .Y(n52) );
  INVX1 U47 ( .A(n37), .Y(n49) );
  MUX2X1 U48 ( .B(n35), .A(n42), .S(n1), .Y(n45) );
  NAND3X1 U49 ( .A(n8), .B(n1), .C(n52), .Y(n43) );
  OAI21X1 U50 ( .A(n29), .B(n41), .C(n27), .Y(n44) );
  OAI21X1 U51 ( .A(n35), .B(n33), .C(n31), .Y(RegDst) );
  AND2X2 U52 ( .A(n39), .B(n4), .Y(n47) );
  AND2X2 U53 ( .A(n47), .B(n46), .Y(writeR7) );
  NAND3X1 U54 ( .A(\opcode<4> ), .B(\opcode<3> ), .C(\opcode<0> ), .Y(n48) );
  NAND3X1 U55 ( .A(\opcode<4> ), .B(n52), .C(\opcode<0> ), .Y(n53) );
endmodule


module writeback ( .nxt_pc({\nxt_pc<15> , \nxt_pc<14> , \nxt_pc<13> , 
        \nxt_pc<12> , \nxt_pc<11> , \nxt_pc<10> , \nxt_pc<9> , \nxt_pc<8> , 
        \nxt_pc<7> , \nxt_pc<6> , \nxt_pc<5> , \nxt_pc<4> , \nxt_pc<3> , 
        \nxt_pc<2> , \nxt_pc<1> , \nxt_pc<0> }), wr_r7, .rd({\rd<2> , \rd<1> , 
        \rd<0> }), .rs({\rs<2> , \rs<1> , \rs<0> }), regdst, memtoreg, slbi, 
        compareS, btr_cntl, .aluOut({\aluOut<15> , \aluOut<14> , \aluOut<13> , 
        \aluOut<12> , \aluOut<11> , \aluOut<10> , \aluOut<9> , \aluOut<8> , 
        \aluOut<7> , \aluOut<6> , \aluOut<5> , \aluOut<4> , \aluOut<3> , 
        \aluOut<2> , \aluOut<1> , \aluOut<0> }), .mem_out({\mem_out<15> , 
        \mem_out<14> , \mem_out<13> , \mem_out<12> , \mem_out<11> , 
        \mem_out<10> , \mem_out<9> , \mem_out<8> , \mem_out<7> , \mem_out<6> , 
        \mem_out<5> , \mem_out<4> , \mem_out<3> , \mem_out<2> , \mem_out<1> , 
        \mem_out<0> }), .alu_out({\alu_out<15> , \alu_out<14> , \alu_out<13> , 
        \alu_out<12> , \alu_out<11> , \alu_out<10> , \alu_out<9> , 
        \alu_out<8> , \alu_out<7> , \alu_out<6> , \alu_out<5> , \alu_out<4> , 
        \alu_out<3> , \alu_out<2> , \alu_out<1> , \alu_out<0> }), .imm({
        \imm<15> , \imm<14> , \imm<13> , \imm<12> , \imm<11> , \imm<10> , 
        \imm<9> , \imm<8> , \imm<7> , \imm<6> , \imm<5> , \imm<4> , \imm<3> , 
        \imm<2> , \imm<1> , \imm<0> }), .writereg({\writereg<2> , 
        \writereg<1> , \writereg<0> }), ofl, zero, N, P, cout, .inst({
        \inst<15> , \inst<14> , \inst<13> , \inst<12> , \inst<11> , \inst<10> , 
        \inst<9> , \inst<8> , \inst<7> , \inst<6> , \inst<5> , \inst<4> , 
        \inst<3> , \inst<2> , \inst<1> , \inst<0> }), ld_imm, .regwritedata({
        \regwritedata<15> , \regwritedata<14> , \regwritedata<13> , 
        \regwritedata<12> , \regwritedata<11> , \regwritedata<10> , 
        \regwritedata<9> , \regwritedata<8> , \regwritedata<7> , 
        \regwritedata<6> , \regwritedata<5> , \regwritedata<4> , 
        \regwritedata<3> , \regwritedata<2> , \regwritedata<1> , 
        \regwritedata<0> }) );
  input \nxt_pc<15> , \nxt_pc<14> , \nxt_pc<13> , \nxt_pc<12> , \nxt_pc<11> ,
         \nxt_pc<10> , \nxt_pc<9> , \nxt_pc<8> , \nxt_pc<7> , \nxt_pc<6> ,
         \nxt_pc<5> , \nxt_pc<4> , \nxt_pc<3> , \nxt_pc<2> , \nxt_pc<1> ,
         \nxt_pc<0> , wr_r7, \rd<2> , \rd<1> , \rd<0> , \rs<2> , \rs<1> ,
         \rs<0> , regdst, memtoreg, slbi, compareS, btr_cntl, \aluOut<15> ,
         \aluOut<14> , \aluOut<13> , \aluOut<12> , \aluOut<11> , \aluOut<10> ,
         \aluOut<9> , \aluOut<8> , \aluOut<7> , \aluOut<6> , \aluOut<5> ,
         \aluOut<4> , \aluOut<3> , \aluOut<2> , \aluOut<1> , \aluOut<0> ,
         \mem_out<15> , \mem_out<14> , \mem_out<13> , \mem_out<12> ,
         \mem_out<11> , \mem_out<10> , \mem_out<9> , \mem_out<8> ,
         \mem_out<7> , \mem_out<6> , \mem_out<5> , \mem_out<4> , \mem_out<3> ,
         \mem_out<2> , \mem_out<1> , \mem_out<0> , \alu_out<15> ,
         \alu_out<14> , \alu_out<13> , \alu_out<12> , \alu_out<11> ,
         \alu_out<10> , \alu_out<9> , \alu_out<8> , \alu_out<7> , \alu_out<6> ,
         \alu_out<5> , \alu_out<4> , \alu_out<3> , \alu_out<2> , \alu_out<1> ,
         \alu_out<0> , \imm<15> , \imm<14> , \imm<13> , \imm<12> , \imm<11> ,
         \imm<10> , \imm<9> , \imm<8> , \imm<7> , \imm<6> , \imm<5> , \imm<4> ,
         \imm<3> , \imm<2> , \imm<1> , \imm<0> , ofl, zero, N, P, cout,
         \inst<15> , \inst<14> , \inst<13> , \inst<12> , \inst<11> ,
         \inst<10> , \inst<9> , \inst<8> , \inst<7> , \inst<6> , \inst<5> ,
         \inst<4> , \inst<3> , \inst<2> , \inst<1> , \inst<0> , ld_imm;
  output \writereg<2> , \writereg<1> , \writereg<0> , \regwritedata<15> ,
         \regwritedata<14> , \regwritedata<13> , \regwritedata<12> ,
         \regwritedata<11> , \regwritedata<10> , \regwritedata<9> ,
         \regwritedata<8> , \regwritedata<7> , \regwritedata<6> ,
         \regwritedata<5> , \regwritedata<4> , \regwritedata<3> ,
         \regwritedata<2> , \regwritedata<1> , \regwritedata<0> ;
  wire   n472, n473, n7, n17, n18, n19, n1, n2, n3, n4, n5, n6, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n307, n308, n309, n310, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471;

  AOI22X1 U23 ( .A(regdst), .B(\rd<2> ), .C(\rs<2> ), .D(n7), .Y(n17) );
  AOI22X1 U24 ( .A(\rd<1> ), .B(regdst), .C(\rs<1> ), .D(n7), .Y(n18) );
  AOI22X1 U25 ( .A(\rd<0> ), .B(regdst), .C(\rs<0> ), .D(n7), .Y(n19) );
  INVX1 U2 ( .A(n362), .Y(n1) );
  BUFX2 U3 ( .A(btr_cntl), .Y(n2) );
  BUFX2 U4 ( .A(btr_cntl), .Y(n3) );
  INVX1 U5 ( .A(n3), .Y(n4) );
  BUFX4 U6 ( .A(btr_cntl), .Y(n360) );
  INVX1 U7 ( .A(\inst<15> ), .Y(n47) );
  INVX1 U8 ( .A(P), .Y(n364) );
  INVX1 U9 ( .A(\mem_out<4> ), .Y(n396) );
  INVX1 U10 ( .A(\mem_out<12> ), .Y(n457) );
  INVX1 U11 ( .A(\nxt_pc<10> ), .Y(n12) );
  INVX1 U12 ( .A(\nxt_pc<12> ), .Y(n37) );
  INVX1 U13 ( .A(\aluOut<3> ), .Y(n455) );
  INVX1 U14 ( .A(\mem_out<13> ), .Y(n461) );
  INVX1 U15 ( .A(\mem_out<14> ), .Y(n465) );
  INVX1 U16 ( .A(\mem_out<15> ), .Y(n469) );
  INVX1 U17 ( .A(\nxt_pc<15> ), .Y(n64) );
  INVX1 U18 ( .A(\aluOut<0> ), .Y(n468) );
  INVX1 U19 ( .A(\aluOut<8> ), .Y(n427) );
  INVX1 U20 ( .A(\inst<14> ), .Y(n49) );
  INVX1 U21 ( .A(\nxt_pc<4> ), .Y(n393) );
  INVX1 U22 ( .A(\imm<5> ), .Y(n404) );
  INVX1 U26 ( .A(\aluOut<14> ), .Y(n371) );
  INVX1 U27 ( .A(\aluOut<13> ), .Y(n379) );
  INVX1 U28 ( .A(\aluOut<6> ), .Y(n430) );
  INVX1 U29 ( .A(\imm<12> ), .Y(n72) );
  INVX1 U30 ( .A(\aluOut<2> ), .Y(n460) );
  INVX1 U31 ( .A(n41), .Y(\regwritedata<15> ) );
  INVX1 U32 ( .A(n440), .Y(n54) );
  INVX1 U33 ( .A(n325), .Y(n38) );
  INVX1 U34 ( .A(n75), .Y(\regwritedata<10> ) );
  OAI21X1 U35 ( .A(n31), .B(n97), .C(n262), .Y(n5) );
  INVX2 U36 ( .A(n4), .Y(n31) );
  INVX1 U37 ( .A(n115), .Y(n6) );
  INVX1 U38 ( .A(n1), .Y(n8) );
  BUFX2 U39 ( .A(n323), .Y(n9) );
  INVX1 U40 ( .A(n339), .Y(n10) );
  NOR3X1 U41 ( .A(n12), .B(n335), .C(n125), .Y(n11) );
  INVX1 U42 ( .A(n334), .Y(n322) );
  INVX1 U43 ( .A(n31), .Y(n13) );
  INVX4 U44 ( .A(n358), .Y(n70) );
  INVX1 U45 ( .A(\inst<13> ), .Y(n48) );
  AND2X2 U46 ( .A(n338), .B(n54), .Y(n14) );
  INVX1 U47 ( .A(n14), .Y(n415) );
  INVX1 U48 ( .A(compareS), .Y(n15) );
  INVX1 U49 ( .A(compareS), .Y(n16) );
  INVX1 U50 ( .A(n338), .Y(n332) );
  INVX1 U51 ( .A(memtoreg), .Y(n338) );
  INVX1 U52 ( .A(n200), .Y(n20) );
  INVX1 U53 ( .A(n200), .Y(n21) );
  INVX1 U54 ( .A(n200), .Y(n22) );
  INVX1 U55 ( .A(n200), .Y(n23) );
  INVX1 U56 ( .A(n429), .Y(n24) );
  INVX1 U57 ( .A(n429), .Y(n25) );
  INVX1 U58 ( .A(n448), .Y(n26) );
  INVX1 U59 ( .A(n448), .Y(n27) );
  INVX1 U60 ( .A(n23), .Y(n28) );
  INVX1 U61 ( .A(n22), .Y(n29) );
  AND2X2 U62 ( .A(\imm<4> ), .B(n65), .Y(n30) );
  NOR2X1 U63 ( .A(n30), .B(n400), .Y(n401) );
  BUFX2 U64 ( .A(compareS), .Y(n361) );
  INVX2 U65 ( .A(n338), .Y(n329) );
  OR2X2 U66 ( .A(n134), .B(n205), .Y(n32) );
  AND2X2 U67 ( .A(n2), .B(n9), .Y(n33) );
  AND2X2 U68 ( .A(n42), .B(n9), .Y(n34) );
  AND2X2 U69 ( .A(n34), .B(n35), .Y(n134) );
  AND2X2 U70 ( .A(n176), .B(n70), .Y(n35) );
  OAI21X1 U71 ( .A(n37), .B(n38), .C(n247), .Y(n36) );
  INVX1 U72 ( .A(n36), .Y(n459) );
  INVX1 U73 ( .A(n88), .Y(n39) );
  INVX1 U74 ( .A(n45), .Y(\regwritedata<5> ) );
  INVX1 U75 ( .A(n359), .Y(n419) );
  OAI21X1 U76 ( .A(n29), .B(n266), .C(n246), .Y(n40) );
  NOR3X1 U77 ( .A(n296), .B(n203), .C(n63), .Y(n41) );
  INVX1 U78 ( .A(n360), .Y(n42) );
  OR2X2 U79 ( .A(n139), .B(n44), .Y(\regwritedata<0> ) );
  INVX1 U80 ( .A(n370), .Y(n44) );
  NOR3X1 U81 ( .A(n40), .B(n255), .C(n293), .Y(n45) );
  INVX1 U82 ( .A(n357), .Y(n65) );
  NOR3X1 U83 ( .A(n47), .B(n48), .C(n49), .Y(n46) );
  INVX1 U84 ( .A(n46), .Y(n365) );
  INVX1 U85 ( .A(n194), .Y(\regwritedata<1> ) );
  AND2X2 U86 ( .A(n167), .B(n180), .Y(n50) );
  OR2X2 U87 ( .A(\inst<12> ), .B(n364), .Y(n269) );
  AND2X2 U88 ( .A(P), .B(\inst<12> ), .Y(n264) );
  INVX1 U89 ( .A(n436), .Y(n51) );
  INVX1 U90 ( .A(n51), .Y(n52) );
  OR2X2 U91 ( .A(n16), .B(n54), .Y(n53) );
  INVX1 U92 ( .A(n53), .Y(n315) );
  INVX1 U93 ( .A(n328), .Y(n55) );
  INVX1 U94 ( .A(n328), .Y(n56) );
  INVX1 U95 ( .A(n56), .Y(n57) );
  INVX1 U96 ( .A(n324), .Y(n58) );
  INVX1 U97 ( .A(n181), .Y(n363) );
  AND2X2 U98 ( .A(cout), .B(\inst<12> ), .Y(n212) );
  INVX1 U99 ( .A(n337), .Y(n328) );
  INVX1 U100 ( .A(n61), .Y(n425) );
  INVX1 U101 ( .A(n89), .Y(n59) );
  INVX1 U102 ( .A(n436), .Y(n60) );
  NOR3X1 U103 ( .A(n178), .B(n62), .C(n188), .Y(n61) );
  INVX1 U104 ( .A(n424), .Y(n62) );
  INVX1 U105 ( .A(wr_r7), .Y(n334) );
  INVX1 U106 ( .A(n351), .Y(\regwritedata<13> ) );
  OAI21X1 U107 ( .A(n64), .B(n38), .C(n252), .Y(n63) );
  INVX1 U108 ( .A(n357), .Y(n470) );
  INVX1 U109 ( .A(wr_r7), .Y(n335) );
  BUFX2 U110 ( .A(ld_imm), .Y(n80) );
  NOR3X1 U111 ( .A(n177), .B(n279), .C(n67), .Y(n66) );
  INVX1 U112 ( .A(n372), .Y(n67) );
  INVX1 U113 ( .A(n102), .Y(n68) );
  INVX1 U114 ( .A(n69), .Y(n456) );
  NOR3X1 U115 ( .A(n93), .B(n321), .C(n326), .Y(n69) );
  AND2X2 U116 ( .A(n87), .B(n207), .Y(n174) );
  OR2X2 U117 ( .A(n318), .B(n460), .Y(n249) );
  BUFX2 U118 ( .A(btr_cntl), .Y(n359) );
  INVX1 U119 ( .A(n358), .Y(n331) );
  OR2X2 U120 ( .A(zero), .B(\inst<11> ), .Y(n267) );
  AND2X2 U121 ( .A(wr_r7), .B(n440), .Y(n297) );
  OAI21X1 U122 ( .A(n72), .B(n357), .C(n248), .Y(n71) );
  INVX1 U123 ( .A(n71), .Y(n458) );
  INVX1 U124 ( .A(n367), .Y(n79) );
  OR2X2 U125 ( .A(n320), .B(n457), .Y(n248) );
  OAI21X1 U126 ( .A(n5), .B(n74), .C(n66), .Y(n73) );
  INVX1 U127 ( .A(n374), .Y(n74) );
  NOR3X1 U128 ( .A(n76), .B(n210), .C(n256), .Y(n75) );
  INVX1 U129 ( .A(n446), .Y(n76) );
  AND2X2 U130 ( .A(n22), .B(n312), .Y(n434) );
  INVX1 U131 ( .A(n77), .Y(n433) );
  NOR3X1 U132 ( .A(n174), .B(n122), .C(n81), .Y(n77) );
  AND2X2 U133 ( .A(n79), .B(n315), .Y(n78) );
  OR2X2 U134 ( .A(compareS), .B(n460), .Y(n286) );
  OR2X2 U135 ( .A(compareS), .B(n393), .Y(n198) );
  OR2X2 U136 ( .A(n243), .B(n361), .Y(n214) );
  AND2X2 U137 ( .A(n361), .B(n440), .Y(n284) );
  OR2X2 U138 ( .A(n6), .B(n428), .Y(n206) );
  OR2X2 U139 ( .A(n358), .B(n360), .Y(n277) );
  AND2X2 U140 ( .A(\imm<10> ), .B(n80), .Y(n226) );
  OR2X2 U141 ( .A(n358), .B(n335), .Y(n257) );
  AND2X2 U142 ( .A(\imm<3> ), .B(n80), .Y(n224) );
  AND2X2 U143 ( .A(n90), .B(n231), .Y(n81) );
  OR2X2 U144 ( .A(n239), .B(n57), .Y(n82) );
  INVX1 U145 ( .A(n82), .Y(n83) );
  OR2X2 U146 ( .A(n197), .B(n85), .Y(\regwritedata<3> ) );
  OR2X2 U147 ( .A(n195), .B(n196), .Y(n85) );
  AND2X2 U148 ( .A(n458), .B(n158), .Y(n86) );
  OR2X2 U149 ( .A(n332), .B(n51), .Y(n429) );
  AND2X2 U150 ( .A(\nxt_pc<9> ), .B(n319), .Y(n87) );
  AND2X2 U151 ( .A(n360), .B(n323), .Y(n88) );
  AND2X2 U152 ( .A(n360), .B(n440), .Y(n89) );
  AND2X2 U153 ( .A(\imm<9> ), .B(n156), .Y(n90) );
  AND2X2 U154 ( .A(n15), .B(n334), .Y(n91) );
  AND2X2 U155 ( .A(\aluOut<11> ), .B(n59), .Y(n92) );
  AND2X2 U156 ( .A(n440), .B(n154), .Y(n93) );
  AND2X2 U157 ( .A(n162), .B(n153), .Y(n94) );
  AND2X2 U158 ( .A(\nxt_pc<0> ), .B(wr_r7), .Y(n95) );
  INVX1 U159 ( .A(n95), .Y(n96) );
  AND2X2 U160 ( .A(\nxt_pc<1> ), .B(wr_r7), .Y(n97) );
  AND2X2 U161 ( .A(\nxt_pc<2> ), .B(n440), .Y(n98) );
  INVX1 U162 ( .A(n98), .Y(n99) );
  AND2X2 U163 ( .A(\imm<2> ), .B(n80), .Y(n100) );
  INVX1 U164 ( .A(n100), .Y(n101) );
  AND2X2 U165 ( .A(n23), .B(n33), .Y(n102) );
  AND2X2 U166 ( .A(\aluOut<4> ), .B(n59), .Y(n103) );
  INVX1 U167 ( .A(n103), .Y(n104) );
  AND2X2 U168 ( .A(n237), .B(n151), .Y(n105) );
  INVX1 U169 ( .A(n105), .Y(\regwritedata<4> ) );
  AND2X2 U170 ( .A(\aluOut<10> ), .B(n3), .Y(n107) );
  INVX1 U171 ( .A(n107), .Y(n108) );
  AND2X2 U172 ( .A(\mem_out<5> ), .B(n329), .Y(n109) );
  INVX1 U173 ( .A(n109), .Y(n110) );
  OR2X2 U174 ( .A(n166), .B(n329), .Y(n111) );
  INVX1 U175 ( .A(n111), .Y(n112) );
  AND2X2 U176 ( .A(n209), .B(n25), .Y(n113) );
  INVX1 U177 ( .A(n113), .Y(n114) );
  AND2X2 U178 ( .A(wr_r7), .B(n42), .Y(n115) );
  AND2X2 U179 ( .A(\nxt_pc<7> ), .B(n191), .Y(n116) );
  INVX1 U180 ( .A(n116), .Y(n117) );
  OR2X2 U181 ( .A(n399), .B(n28), .Y(n118) );
  INVX1 U182 ( .A(n118), .Y(n119) );
  AND2X2 U183 ( .A(n160), .B(n152), .Y(n120) );
  INVX1 U184 ( .A(n120), .Y(\regwritedata<7> ) );
  AND2X2 U185 ( .A(\mem_out<9> ), .B(n356), .Y(n122) );
  AND2X2 U186 ( .A(n319), .B(n211), .Y(n123) );
  INVX1 U187 ( .A(n123), .Y(n124) );
  OR2X2 U188 ( .A(n332), .B(n360), .Y(n125) );
  INVX1 U189 ( .A(n125), .Y(n126) );
  AND2X2 U190 ( .A(\mem_out<11> ), .B(n356), .Y(n127) );
  INVX1 U191 ( .A(n127), .Y(n128) );
  AND2X2 U192 ( .A(\nxt_pc<14> ), .B(n325), .Y(n129) );
  INVX1 U193 ( .A(n129), .Y(n130) );
  AND2X2 U194 ( .A(\aluOut<14> ), .B(n345), .Y(n131) );
  INVX1 U195 ( .A(n131), .Y(n132) );
  BUFX2 U196 ( .A(n463), .Y(n133) );
  AND2X2 U197 ( .A(n356), .B(\mem_out<7> ), .Y(n135) );
  INVX1 U198 ( .A(n135), .Y(n136) );
  OR2X2 U199 ( .A(n429), .B(n58), .Y(n137) );
  INVX1 U200 ( .A(n137), .Y(n138) );
  OR2X2 U201 ( .A(n32), .B(n330), .Y(n139) );
  AND2X2 U202 ( .A(n319), .B(n78), .Y(n140) );
  INVX1 U203 ( .A(n140), .Y(n141) );
  OR2X2 U204 ( .A(n99), .B(compareS), .Y(n142) );
  INVX1 U205 ( .A(n142), .Y(n143) );
  AND2X2 U206 ( .A(\imm<7> ), .B(n470), .Y(n144) );
  INVX1 U207 ( .A(n144), .Y(n145) );
  BUFX2 U208 ( .A(n376), .Y(n146) );
  BUFX2 U209 ( .A(n395), .Y(n147) );
  BUFX2 U210 ( .A(n426), .Y(n148) );
  AND2X2 U211 ( .A(n202), .B(n23), .Y(n149) );
  INVX1 U212 ( .A(n149), .Y(n150) );
  BUFX2 U213 ( .A(n401), .Y(n151) );
  BUFX2 U214 ( .A(n423), .Y(n152) );
  BUFX2 U215 ( .A(n462), .Y(n153) );
  INVX1 U216 ( .A(n91), .Y(n154) );
  AND2X2 U217 ( .A(n440), .B(n331), .Y(n155) );
  INVX1 U218 ( .A(n155), .Y(n156) );
  AND2X2 U219 ( .A(\aluOut<12> ), .B(n344), .Y(n157) );
  INVX1 U220 ( .A(n157), .Y(n158) );
  OR2X2 U221 ( .A(n164), .B(n420), .Y(n159) );
  INVX1 U222 ( .A(n159), .Y(n160) );
  AND2X2 U223 ( .A(\aluOut<13> ), .B(n345), .Y(n161) );
  INVX1 U224 ( .A(n161), .Y(n162) );
  AND2X2 U225 ( .A(n145), .B(n136), .Y(n163) );
  INVX1 U226 ( .A(n163), .Y(n164) );
  AND2X2 U227 ( .A(n322), .B(n229), .Y(n165) );
  INVX1 U228 ( .A(n165), .Y(n166) );
  AND2X2 U229 ( .A(\aluOut<0> ), .B(n59), .Y(n167) );
  AND2X2 U230 ( .A(n322), .B(n143), .Y(n168) );
  INVX1 U231 ( .A(n168), .Y(n169) );
  BUFX2 U232 ( .A(n453), .Y(n170) );
  AND2X2 U233 ( .A(n235), .B(n141), .Y(n171) );
  INVX1 U234 ( .A(n171), .Y(n172) );
  BUFX2 U235 ( .A(n381), .Y(n173) );
  OR2X2 U236 ( .A(n96), .B(n362), .Y(n175) );
  INVX1 U237 ( .A(n175), .Y(n176) );
  AND2X2 U238 ( .A(\imm<1> ), .B(n80), .Y(n177) );
  AND2X2 U239 ( .A(\mem_out<8> ), .B(n356), .Y(n178) );
  BUFX2 U240 ( .A(n473), .Y(\regwritedata<2> ) );
  OR2X2 U241 ( .A(n91), .B(slbi), .Y(n180) );
  INVX1 U242 ( .A(n180), .Y(n181) );
  OR2X2 U243 ( .A(n169), .B(n358), .Y(n182) );
  INVX1 U244 ( .A(n182), .Y(n183) );
  AND2X2 U245 ( .A(n92), .B(n363), .Y(n184) );
  INVX1 U246 ( .A(n184), .Y(n185) );
  OR2X2 U247 ( .A(n379), .B(n316), .Y(n186) );
  INVX1 U248 ( .A(n186), .Y(n187) );
  AND2X2 U249 ( .A(\imm<8> ), .B(n65), .Y(n188) );
  OR2X2 U250 ( .A(slbi), .B(compareS), .Y(n189) );
  INVX1 U251 ( .A(n189), .Y(n190) );
  INVX1 U252 ( .A(n189), .Y(n191) );
  AND2X2 U253 ( .A(n86), .B(n459), .Y(n192) );
  INVX1 U254 ( .A(n192), .Y(\regwritedata<12> ) );
  BUFX2 U255 ( .A(n353), .Y(n194) );
  INVX1 U256 ( .A(n392), .Y(n195) );
  INVX1 U257 ( .A(n391), .Y(n196) );
  INVX1 U258 ( .A(n390), .Y(n197) );
  INVX1 U259 ( .A(n198), .Y(n199) );
  INVX1 U260 ( .A(n320), .Y(n410) );
  OR2X2 U261 ( .A(n328), .B(n60), .Y(n200) );
  OR2X2 U262 ( .A(n39), .B(n430), .Y(n201) );
  INVX1 U263 ( .A(n201), .Y(n202) );
  AND2X2 U264 ( .A(\aluOut<15> ), .B(n345), .Y(n203) );
  OR2X2 U265 ( .A(n233), .B(n461), .Y(n204) );
  INVX1 U266 ( .A(n369), .Y(n205) );
  INVX1 U267 ( .A(n206), .Y(n207) );
  OR2X2 U268 ( .A(n245), .B(n2), .Y(n208) );
  INVX1 U269 ( .A(n208), .Y(n209) );
  INVX1 U270 ( .A(n445), .Y(n210) );
  INVX1 U271 ( .A(n190), .Y(n428) );
  INVX1 U272 ( .A(regdst), .Y(n7) );
  INVX1 U273 ( .A(n89), .Y(n211) );
  INVX1 U274 ( .A(n212), .Y(n213) );
  INVX1 U275 ( .A(n214), .Y(n215) );
  INVX1 U276 ( .A(n412), .Y(n216) );
  INVX1 U277 ( .A(n216), .Y(n217) );
  INVX1 U278 ( .A(n366), .Y(n218) );
  INVX1 U279 ( .A(n218), .Y(n219) );
  INVX1 U280 ( .A(n447), .Y(n220) );
  INVX1 U281 ( .A(n220), .Y(n221) );
  INVX1 U282 ( .A(n464), .Y(n222) );
  INVX1 U283 ( .A(n222), .Y(n223) );
  INVX1 U284 ( .A(n224), .Y(n225) );
  INVX1 U285 ( .A(n226), .Y(n227) );
  OR2X2 U286 ( .A(n241), .B(compareS), .Y(n228) );
  INVX1 U287 ( .A(n228), .Y(n229) );
  INVX1 U288 ( .A(n233), .Y(n230) );
  INVX1 U289 ( .A(n230), .Y(n231) );
  AND2X2 U290 ( .A(n52), .B(n362), .Y(n232) );
  INVX1 U291 ( .A(n232), .Y(n233) );
  INVX1 U292 ( .A(n368), .Y(n234) );
  INVX1 U293 ( .A(n234), .Y(n235) );
  INVX1 U294 ( .A(n402), .Y(n236) );
  INVX1 U295 ( .A(n236), .Y(n237) );
  AND2X1 U296 ( .A(\imm<0> ), .B(slbi), .Y(n238) );
  INVX1 U297 ( .A(n238), .Y(n239) );
  AND2X2 U298 ( .A(\nxt_pc<5> ), .B(n440), .Y(n240) );
  INVX1 U299 ( .A(n240), .Y(n241) );
  AND2X1 U300 ( .A(\aluOut<9> ), .B(n440), .Y(n242) );
  INVX1 U301 ( .A(n242), .Y(n243) );
  AND2X2 U302 ( .A(\nxt_pc<6> ), .B(wr_r7), .Y(n244) );
  INVX1 U303 ( .A(n244), .Y(n245) );
  OR2X2 U304 ( .A(n110), .B(n80), .Y(n246) );
  OR2X2 U305 ( .A(n68), .B(n455), .Y(n247) );
  INVX1 U306 ( .A(n249), .Y(n250) );
  INVX1 U307 ( .A(n204), .Y(n251) );
  OR2X2 U308 ( .A(n318), .B(n468), .Y(n252) );
  OR2X2 U309 ( .A(n233), .B(n469), .Y(n253) );
  INVX1 U310 ( .A(n253), .Y(n254) );
  INVX1 U311 ( .A(n407), .Y(n255) );
  INVX1 U312 ( .A(n444), .Y(n256) );
  INVX1 U313 ( .A(n257), .Y(n258) );
  BUFX2 U314 ( .A(n19), .Y(n259) );
  INVX1 U315 ( .A(n259), .Y(\writereg<0> ) );
  BUFX2 U316 ( .A(n18), .Y(n260) );
  INVX1 U317 ( .A(n260), .Y(\writereg<1> ) );
  BUFX2 U318 ( .A(n17), .Y(n261) );
  INVX1 U319 ( .A(n261), .Y(\writereg<2> ) );
  AND2X2 U320 ( .A(n191), .B(n55), .Y(n262) );
  INVX1 U321 ( .A(n262), .Y(n263) );
  INVX1 U322 ( .A(n263), .Y(n450) );
  INVX1 U323 ( .A(n264), .Y(n265) );
  OR2X2 U324 ( .A(n108), .B(n428), .Y(n266) );
  INVX1 U325 ( .A(n267), .Y(n268) );
  INVX1 U326 ( .A(n269), .Y(n270) );
  AND2X1 U327 ( .A(\imm<2> ), .B(slbi), .Y(n271) );
  INVX1 U328 ( .A(n271), .Y(n272) );
  AND2X1 U329 ( .A(\imm<3> ), .B(slbi), .Y(n273) );
  INVX1 U330 ( .A(n273), .Y(n274) );
  AND2X1 U331 ( .A(\imm<10> ), .B(slbi), .Y(n275) );
  INVX1 U332 ( .A(n275), .Y(n276) );
  INVX1 U333 ( .A(n277), .Y(n278) );
  INVX1 U334 ( .A(n373), .Y(n279) );
  INVX1 U335 ( .A(n382), .Y(n280) );
  INVX1 U336 ( .A(n280), .Y(n281) );
  INVX1 U337 ( .A(n451), .Y(n282) );
  INVX1 U338 ( .A(n282), .Y(n283) );
  INVX1 U339 ( .A(n284), .Y(n285) );
  INVX1 U340 ( .A(n286), .Y(n287) );
  BUFX2 U341 ( .A(n431), .Y(n288) );
  AND2X2 U342 ( .A(\inst<11> ), .B(n213), .Y(n289) );
  INVX1 U343 ( .A(n289), .Y(n290) );
  INVX1 U344 ( .A(n405), .Y(n291) );
  INVX1 U345 ( .A(n291), .Y(n292) );
  INVX1 U346 ( .A(n406), .Y(n293) );
  INVX1 U347 ( .A(n467), .Y(n294) );
  INVX1 U348 ( .A(n294), .Y(n295) );
  INVX1 U349 ( .A(n471), .Y(n296) );
  INVX1 U350 ( .A(n297), .Y(n298) );
  AND2X1 U351 ( .A(\aluOut<12> ), .B(n440), .Y(n299) );
  INVX1 U352 ( .A(n299), .Y(n300) );
  AND2X1 U353 ( .A(\aluOut<5> ), .B(n440), .Y(n301) );
  INVX1 U354 ( .A(n301), .Y(n302) );
  INVX1 U355 ( .A(n11), .Y(n303) );
  INVX1 U356 ( .A(n232), .Y(n304) );
  INVX1 U357 ( .A(n472), .Y(n305) );
  INVX1 U358 ( .A(n305), .Y(\regwritedata<14> ) );
  INVX1 U359 ( .A(n308), .Y(n307) );
  AND2X1 U360 ( .A(\aluOut<6> ), .B(slbi), .Y(n308) );
  INVX1 U361 ( .A(n115), .Y(n309) );
  INVX1 U362 ( .A(n297), .Y(n310) );
  INVX1 U363 ( .A(n89), .Y(n312) );
  INVX1 U364 ( .A(n53), .Y(n313) );
  INVX1 U365 ( .A(n313), .Y(n314) );
  INVX1 U366 ( .A(n324), .Y(n316) );
  INVX1 U367 ( .A(n88), .Y(n317) );
  INVX1 U368 ( .A(n102), .Y(n318) );
  INVX1 U369 ( .A(n200), .Y(n319) );
  INVX1 U370 ( .A(n232), .Y(n320) );
  AND2X2 U371 ( .A(n3), .B(n440), .Y(n321) );
  INVX1 U372 ( .A(memtoreg), .Y(n337) );
  INVX1 U373 ( .A(n191), .Y(n437) );
  AND2X2 U374 ( .A(n440), .B(n336), .Y(n323) );
  AND2X2 U375 ( .A(n359), .B(n323), .Y(n324) );
  AND2X2 U376 ( .A(n333), .B(n450), .Y(n325) );
  INVX1 U377 ( .A(n342), .Y(n326) );
  INVX1 U378 ( .A(n414), .Y(n327) );
  INVX1 U379 ( .A(n2), .Y(n441) );
  AND2X2 U380 ( .A(n138), .B(\aluOut<15> ), .Y(n330) );
  INVX1 U381 ( .A(n337), .Y(n362) );
  NOR3X1 U382 ( .A(n3), .B(n358), .C(n335), .Y(n333) );
  INVX1 U383 ( .A(n375), .Y(n354) );
  INVX1 U384 ( .A(ld_imm), .Y(n436) );
  INVX1 U385 ( .A(compareS), .Y(n336) );
  INVX1 U386 ( .A(n414), .Y(n339) );
  INVX1 U387 ( .A(n339), .Y(n340) );
  INVX1 U388 ( .A(n342), .Y(n341) );
  INVX1 U389 ( .A(n414), .Y(n342) );
  INVX1 U390 ( .A(n345), .Y(n343) );
  INVX1 U391 ( .A(n456), .Y(n344) );
  INVX1 U392 ( .A(n180), .Y(n399) );
  INVX1 U393 ( .A(n456), .Y(n345) );
  OR2X2 U394 ( .A(n329), .B(n349), .Y(n346) );
  AND2X2 U395 ( .A(n346), .B(n347), .Y(n452) );
  OR2X2 U396 ( .A(n70), .B(n348), .Y(n347) );
  INVX1 U397 ( .A(\imm<11> ), .Y(n348) );
  OR2X2 U398 ( .A(n440), .B(n348), .Y(n349) );
  AND2X2 U399 ( .A(n133), .B(n94), .Y(n351) );
  INVX1 U400 ( .A(n377), .Y(n350) );
  OR2X2 U401 ( .A(n350), .B(n10), .Y(n383) );
  INVX1 U402 ( .A(n318), .Y(n398) );
  AOI21X1 U403 ( .A(n355), .B(n354), .C(n73), .Y(n353) );
  AND2X2 U404 ( .A(n312), .B(n25), .Y(n355) );
  INVX1 U405 ( .A(n304), .Y(n356) );
  AND2X2 U406 ( .A(n52), .B(n415), .Y(n357) );
  INVX8 U407 ( .A(slbi), .Y(n440) );
  BUFX4 U408 ( .A(ld_imm), .Y(n358) );
  OR2X2 U409 ( .A(n332), .B(n51), .Y(n448) );
  NAND3X1 U410 ( .A(\mem_out<0> ), .B(n329), .C(n70), .Y(n368) );
  AOI21X1 U411 ( .A(n268), .B(n265), .C(n365), .Y(n366) );
  OAI21X1 U412 ( .A(n270), .B(n290), .C(n219), .Y(n367) );
  AOI21X1 U413 ( .A(n20), .B(n50), .C(n172), .Y(n370) );
  AOI21X1 U414 ( .A(\imm<0> ), .B(n80), .C(n83), .Y(n369) );
  NAND3X1 U415 ( .A(\aluOut<1> ), .B(n285), .C(n298), .Y(n375) );
  AOI21X1 U416 ( .A(n371), .B(n31), .C(n358), .Y(n374) );
  NAND3X1 U417 ( .A(\imm<1> ), .B(slbi), .C(n55), .Y(n373) );
  NAND3X1 U418 ( .A(n329), .B(n331), .C(\mem_out<1> ), .Y(n372) );
  NAND3X1 U419 ( .A(n335), .B(n287), .C(n419), .Y(n376) );
  OAI21X1 U420 ( .A(n440), .B(n460), .C(n146), .Y(n377) );
  OAI21X1 U421 ( .A(n272), .B(n8), .C(n101), .Y(n378) );
  AOI21X1 U422 ( .A(n183), .B(n126), .C(n378), .Y(n382) );
  AND2X2 U423 ( .A(\mem_out<2> ), .B(n329), .Y(n380) );
  AOI22X1 U424 ( .A(n70), .B(n380), .C(n20), .D(n187), .Y(n381) );
  NAND3X1 U425 ( .A(n383), .B(n281), .C(n173), .Y(n473) );
  NOR3X1 U426 ( .A(n2), .B(n428), .C(n335), .Y(n386) );
  AND2X2 U427 ( .A(n21), .B(\nxt_pc<3> ), .Y(n385) );
  OAI21X1 U428 ( .A(n274), .B(n8), .C(n225), .Y(n384) );
  AOI21X1 U429 ( .A(n386), .B(n385), .C(n384), .Y(n392) );
  AND2X2 U430 ( .A(\mem_out<3> ), .B(n329), .Y(n388) );
  NOR3X1 U431 ( .A(n361), .B(n300), .C(n441), .Y(n387) );
  AOI22X1 U432 ( .A(n70), .B(n388), .C(n26), .D(n387), .Y(n391) );
  AND2X2 U433 ( .A(n312), .B(\aluOut<3> ), .Y(n389) );
  NAND3X1 U434 ( .A(n389), .B(n22), .C(n363), .Y(n390) );
  NOR3X1 U435 ( .A(n31), .B(n8), .C(slbi), .Y(n394) );
  NAND3X1 U436 ( .A(n258), .B(n199), .C(n394), .Y(n395) );
  OAI21X1 U437 ( .A(n231), .B(n396), .C(n147), .Y(n397) );
  AOI21X1 U438 ( .A(\aluOut<11> ), .B(n398), .C(n397), .Y(n402) );
  NOR3X1 U439 ( .A(n399), .B(n104), .C(n341), .Y(n400) );
  AND2X2 U440 ( .A(n24), .B(n211), .Y(n403) );
  NAND3X1 U441 ( .A(\aluOut<5> ), .B(n363), .C(n403), .Y(n407) );
  AOI21X1 U442 ( .A(n440), .B(n70), .C(n404), .Y(n405) );
  AOI22X1 U443 ( .A(n278), .B(n112), .C(n320), .D(n292), .Y(n406) );
  OR2X2 U444 ( .A(n358), .B(n57), .Y(n414) );
  OR2X2 U445 ( .A(n361), .B(n430), .Y(n408) );
  OAI21X1 U446 ( .A(n408), .B(n322), .C(n307), .Y(n409) );
  OAI21X1 U447 ( .A(n308), .B(n13), .C(n409), .Y(n413) );
  AND2X2 U448 ( .A(n215), .B(n31), .Y(n411) );
  AOI22X1 U449 ( .A(n21), .B(n411), .C(\mem_out<6> ), .D(n410), .Y(n412) );
  OAI21X1 U450 ( .A(n29), .B(n413), .C(n217), .Y(n418) );
  OAI21X1 U451 ( .A(n14), .B(n80), .C(\imm<6> ), .Y(n416) );
  OAI21X1 U452 ( .A(n428), .B(n114), .C(n416), .Y(n417) );
  OR2X2 U453 ( .A(n417), .B(n418), .Y(\regwritedata<6> ) );
  NOR3X1 U454 ( .A(n341), .B(n309), .C(n117), .Y(n420) );
  AND2X2 U455 ( .A(n211), .B(\aluOut<7> ), .Y(n422) );
  NOR3X1 U456 ( .A(n317), .B(n427), .C(n340), .Y(n421) );
  AOI21X1 U457 ( .A(n422), .B(n119), .C(n421), .Y(n423) );
  NOR3X1 U458 ( .A(n360), .B(n358), .C(n335), .Y(n449) );
  NAND3X1 U459 ( .A(n33), .B(n27), .C(\aluOut<7> ), .Y(n424) );
  AOI21X1 U460 ( .A(\nxt_pc<8> ), .B(n325), .C(n425), .Y(n426) );
  OAI21X1 U461 ( .A(n343), .B(n427), .C(n148), .Y(\regwritedata<8> ) );
  NAND3X1 U462 ( .A(\aluOut<9> ), .B(n314), .C(n310), .Y(n431) );
  OAI21X1 U463 ( .A(n124), .B(n288), .C(n150), .Y(n432) );
  OR2X2 U464 ( .A(n433), .B(n432), .Y(\regwritedata<9> ) );
  AND2X2 U465 ( .A(\aluOut<10> ), .B(n314), .Y(n435) );
  NAND3X1 U466 ( .A(n310), .B(n435), .C(n434), .Y(n446) );
  AND2X2 U467 ( .A(n8), .B(n70), .Y(n439) );
  NOR3X1 U468 ( .A(n80), .B(n437), .C(n303), .Y(n438) );
  AOI21X1 U469 ( .A(n439), .B(\mem_out<10> ), .C(n438), .Y(n445) );
  NOR3X1 U470 ( .A(n441), .B(n302), .C(n361), .Y(n443) );
  OAI21X1 U471 ( .A(n276), .B(n8), .C(n227), .Y(n442) );
  AOI21X1 U472 ( .A(n24), .B(n443), .C(n442), .Y(n444) );
  NAND3X1 U473 ( .A(n33), .B(n20), .C(\aluOut<4> ), .Y(n447) );
  OAI21X1 U474 ( .A(n185), .B(n29), .C(n221), .Y(n454) );
  NAND3X1 U475 ( .A(\nxt_pc<11> ), .B(n450), .C(n449), .Y(n451) );
  NAND3X1 U476 ( .A(n128), .B(n283), .C(n452), .Y(n453) );
  OR2X2 U477 ( .A(n454), .B(n170), .Y(\regwritedata<11> ) );
  AOI21X1 U478 ( .A(\nxt_pc<13> ), .B(n325), .C(n250), .Y(n463) );
  AOI21X1 U479 ( .A(\imm<13> ), .B(n65), .C(n251), .Y(n462) );
  NAND3X1 U480 ( .A(n33), .B(n327), .C(\aluOut<1> ), .Y(n464) );
  OAI21X1 U481 ( .A(n320), .B(n465), .C(n223), .Y(n466) );
  AOI21X1 U482 ( .A(\imm<14> ), .B(n65), .C(n466), .Y(n467) );
  NAND3X1 U483 ( .A(n130), .B(n132), .C(n295), .Y(n472) );
  AOI21X1 U484 ( .A(\imm<15> ), .B(n65), .C(n254), .Y(n471) );
endmodule


module Harzard ( .ID_rs({\ID_rs<2> , \ID_rs<1> , \ID_rs<0> }), .ID_rt({
        \ID_rt<2> , \ID_rt<1> , \ID_rt<0> }), .EX_rd({\EX_rd<2> , \EX_rd<1> , 
        \EX_rd<0> }), .MEM_rd({\MEM_rd<2> , \MEM_rd<1> , \MEM_rd<0> }), 
        ID_rs_v, ID_rt_v, EX_rd_v, MEM_rd_v, .EX_inst({\EX_inst<15> , 
        \EX_inst<14> , \EX_inst<13> , \EX_inst<12> , \EX_inst<11> , 
        \EX_inst<10> , \EX_inst<9> , \EX_inst<8> , \EX_inst<7> , \EX_inst<6> , 
        \EX_inst<5> , \EX_inst<4> , \EX_inst<3> , \EX_inst<2> , \EX_inst<1> , 
        \EX_inst<0> }), .MEM_inst({\MEM_inst<15> , \MEM_inst<14> , 
        \MEM_inst<13> , \MEM_inst<12> , \MEM_inst<11> , \MEM_inst<10> , 
        \MEM_inst<9> , \MEM_inst<8> , \MEM_inst<7> , \MEM_inst<6> , 
        \MEM_inst<5> , \MEM_inst<4> , \MEM_inst<3> , \MEM_inst<2> , 
        \MEM_inst<1> , \MEM_inst<0> }), fow_EXID_rs, fow_EXID_rt, fow_MEMID_rs, 
        fow_MEMID_rt, memStall, memDone, memwrite, memread, stall, 
        instMemStall, instMemDone, instMemDone_q, clk, rst );
  input \ID_rs<2> , \ID_rs<1> , \ID_rs<0> , \ID_rt<2> , \ID_rt<1> , \ID_rt<0> ,
         \EX_rd<2> , \EX_rd<1> , \EX_rd<0> , \MEM_rd<2> , \MEM_rd<1> ,
         \MEM_rd<0> , ID_rs_v, ID_rt_v, EX_rd_v, MEM_rd_v, \EX_inst<15> ,
         \EX_inst<14> , \EX_inst<13> , \EX_inst<12> , \EX_inst<11> ,
         \EX_inst<10> , \EX_inst<9> , \EX_inst<8> , \EX_inst<7> , \EX_inst<6> ,
         \EX_inst<5> , \EX_inst<4> , \EX_inst<3> , \EX_inst<2> , \EX_inst<1> ,
         \EX_inst<0> , \MEM_inst<15> , \MEM_inst<14> , \MEM_inst<13> ,
         \MEM_inst<12> , \MEM_inst<11> , \MEM_inst<10> , \MEM_inst<9> ,
         \MEM_inst<8> , \MEM_inst<7> , \MEM_inst<6> , \MEM_inst<5> ,
         \MEM_inst<4> , \MEM_inst<3> , \MEM_inst<2> , \MEM_inst<1> ,
         \MEM_inst<0> , memStall, memDone, memwrite, memread, instMemStall,
         instMemDone, instMemDone_q, clk, rst;
  output fow_EXID_rs, fow_EXID_rt, fow_MEMID_rs, fow_MEMID_rt, stall;
  wire   n1, n2, n3, n4, n5, n7, n8, n9, n10, n11, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n6, n12, n28, n29,
         n30, n31, n32, n33, n34;

  dff_162 stallq ( .q(), .d(1'b0), .clk(clk), .rst(rst) );
  dff_161 memDoneq ( .q(), .d(memDone), .clk(clk), .rst(rst) );
  dff_160 stallst ( .q(), .d(1'b0), .clk(clk), .rst(rst) );
  OAI21X1 U5 ( .A(instMemDone_q), .B(instMemDone), .C(n4), .Y(stall) );
  OAI21X1 U6 ( .A(memread), .B(memwrite), .C(n3), .Y(n4) );
  NOR3X1 U7 ( .A(n29), .B(n2), .C(n33), .Y(fow_MEMID_rt) );
  NAND3X1 U9 ( .A(n8), .B(n9), .C(n10), .Y(n5) );
  XNOR2X1 U10 ( .A(\ID_rt<1> ), .B(\MEM_rd<1> ), .Y(n10) );
  XNOR2X1 U11 ( .A(\ID_rt<0> ), .B(\MEM_rd<0> ), .Y(n9) );
  XNOR2X1 U12 ( .A(\ID_rt<2> ), .B(\MEM_rd<2> ), .Y(n8) );
  NOR3X1 U13 ( .A(n28), .B(n1), .C(n31), .Y(fow_MEMID_rs) );
  NAND3X1 U15 ( .A(n13), .B(n14), .C(n15), .Y(n7) );
  XNOR2X1 U16 ( .A(\MEM_rd<2> ), .B(\EX_rd<2> ), .Y(n16) );
  XNOR2X1 U17 ( .A(\EX_rd<1> ), .B(\MEM_rd<1> ), .Y(n14) );
  XNOR2X1 U18 ( .A(\EX_rd<0> ), .B(\MEM_rd<0> ), .Y(n13) );
  NAND3X1 U19 ( .A(n17), .B(n18), .C(n19), .Y(n11) );
  XNOR2X1 U20 ( .A(\ID_rs<1> ), .B(\MEM_rd<1> ), .Y(n19) );
  XNOR2X1 U21 ( .A(\ID_rs<0> ), .B(\MEM_rd<0> ), .Y(n18) );
  XNOR2X1 U22 ( .A(\ID_rs<2> ), .B(\MEM_rd<2> ), .Y(n17) );
  NOR3X1 U23 ( .A(n12), .B(n21), .C(n22), .Y(fow_EXID_rt) );
  XOR2X1 U24 ( .A(\ID_rt<0> ), .B(\EX_rd<0> ), .Y(n22) );
  XOR2X1 U25 ( .A(\ID_rt<1> ), .B(\EX_rd<1> ), .Y(n21) );
  NAND3X1 U26 ( .A(ID_rt_v), .B(EX_rd_v), .C(n23), .Y(n20) );
  XNOR2X1 U27 ( .A(\EX_rd<2> ), .B(\ID_rt<2> ), .Y(n23) );
  NOR3X1 U28 ( .A(n6), .B(n25), .C(n26), .Y(fow_EXID_rs) );
  XOR2X1 U29 ( .A(\ID_rs<0> ), .B(\EX_rd<0> ), .Y(n26) );
  XOR2X1 U30 ( .A(\ID_rs<1> ), .B(\EX_rd<1> ), .Y(n25) );
  NAND3X1 U31 ( .A(ID_rs_v), .B(EX_rd_v), .C(n27), .Y(n24) );
  XNOR2X1 U32 ( .A(\EX_rd<2> ), .B(\ID_rs<2> ), .Y(n27) );
  INVX1 U1 ( .A(memDone), .Y(n3) );
  INVX1 U2 ( .A(ID_rs_v), .Y(n1) );
  INVX1 U3 ( .A(MEM_rd_v), .Y(n2) );
  AND2X1 U4 ( .A(EX_rd_v), .B(n16), .Y(n15) );
  BUFX2 U8 ( .A(n24), .Y(n6) );
  BUFX2 U14 ( .A(n20), .Y(n12) );
  BUFX2 U33 ( .A(n11), .Y(n28) );
  BUFX2 U34 ( .A(n5), .Y(n29) );
  AND2X1 U35 ( .A(MEM_rd_v), .B(n34), .Y(n30) );
  INVX1 U36 ( .A(n30), .Y(n31) );
  AND2X1 U37 ( .A(ID_rt_v), .B(n34), .Y(n32) );
  INVX1 U38 ( .A(n32), .Y(n33) );
  BUFX2 U39 ( .A(n7), .Y(n34) );
endmodule


module proc ( err, clk, rst );
  input clk, rst;
  output err;
  wire   stall, jump_IF, jump_ID, br_ctl, pc_en, IcacheErr, DcacheErr,
         rf_bypass_err, instMemDone_q, instMemDone, instMemDone_d,
         \instIF_q<15> , \instIF_q<14> , \instIF_q<13> , \instIF_q<12> ,
         \instIF_q<11> , \instIF_q<10> , \instIF_q<9> , \instIF_q<8> ,
         \instIF_q<7> , \instIF_q<6> , \instIF_q<5> , \instIF_q<4> ,
         \instIF_q<3> , \instIF_q<2> , \instIF_q<1> , \instIF_q<0> , jump_EX,
         \instIF_normal<15> , \instIF_normal<14> , \instIF_normal<13> ,
         \instIF_normal<12> , \instIF_normal<11> , \instIF_normal<10> ,
         \instIF_normal<9> , \instIF_normal<8> , \instIF_normal<7> ,
         \instIF_normal<6> , \instIF_normal<5> , \instIF_normal<4> ,
         \instIF_normal<3> , \instIF_normal<2> , \instIF_normal<1> ,
         \instIF_normal<0> , branch_if, \pc_inc_two<15> , \pc_inc_two<14> ,
         \pc_inc_two<13> , \pc_inc_two<12> , \pc_inc_two<11> ,
         \pc_inc_two<10> , \pc_inc_two<9> , \pc_inc_two<8> , \pc_inc_two<7> ,
         \pc_inc_two<6> , \pc_inc_two<5> , \pc_inc_two<4> , \pc_inc_two<3> ,
         \pc_inc_two<2> , \pc_inc_two<1> , \pc_inc_two<0> , \addr<15> ,
         \addr<14> , \addr<13> , \addr<12> , \addr<11> , \addr<10> , \addr<9> ,
         \addr<8> , \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> ,
         \addr<2> , \addr<1> , \addr<0> , branch_ex,
         \forwarded_read1dataEX<15> , \forwarded_read1dataEX<13> ,
         \forwarded_read1dataEX<12> , \forwarded_read1dataEX<9> ,
         \forwarded_read1dataEX<8> , \forwarded_read1dataEX<5> , \pc_nx<15> ,
         \pc_nx<14> , \pc_nx<13> , \pc_nx<12> , \pc_nx<11> , \pc_nx<10> ,
         \pc_nx<9> , \pc_nx<8> , \pc_nx<7> , \pc_nx<6> , \pc_nx<5> ,
         \pc_nx<4> , \pc_nx<3> , \pc_nx<2> , \pc_nx<1> , \pc_nx<0> ,
         \instEX_normal<15> , \instEX_normal<14> , \instEX_normal<13> ,
         \instEX_normal<12> , \instEX_normal<11> , \instEX_normal<10> ,
         \instEX_normal<9> , \instEX_normal<8> , \instEX_normal<7> ,
         \instEX_normal<6> , \instEX_normal<5> , \instEX_normal<4> ,
         \instEX_normal<3> , \instEX_normal<2> , \instEX_normal<1> ,
         \instEX_normal<0> , instMemStall, _3_net_, haltMEM, \wr_instIF<15> ,
         \wr_instIF<14> , \wr_instIF<13> , \wr_instIF<12> , \wr_instIF<11> ,
         \wr_instIF<10> , \wr_instIF<9> , \wr_instIF<8> , \wr_instIF<7> ,
         \wr_instIF<6> , \wr_instIF<5> , \wr_instIF<4> , \wr_instIF<3> ,
         \wr_instIF<2> , \wr_instIF<1> , \wr_instIF<0> , \instID<15> ,
         \instID<14> , \instID<13> , \instID<12> , \instID<11> , \instID<10> ,
         \instID<9> , \instID<8> , \instID<7> , \instID<6> , \instID<5> ,
         \instID<4> , \instID<3> , \instID<2> , \instID<1> , \instID<0> ,
         \nx_pcID<15> , \nx_pcID<14> , \nx_pcID<13> , \nx_pcID<12> ,
         \nx_pcID<11> , \nx_pcID<10> , \nx_pcID<9> , \nx_pcID<8> ,
         \nx_pcID<7> , \nx_pcID<6> , \nx_pcID<5> , \nx_pcID<4> , \nx_pcID<3> ,
         \nx_pcID<2> , \nx_pcID<1> , \nx_pcID<0> , \pc_inc_two_ID<15> ,
         \pc_inc_two_ID<14> , \pc_inc_two_ID<13> , \pc_inc_two_ID<12> ,
         \pc_inc_two_ID<11> , \pc_inc_two_ID<10> , \pc_inc_two_ID<9> ,
         \pc_inc_two_ID<8> , \pc_inc_two_ID<7> , \pc_inc_two_ID<6> ,
         \pc_inc_two_ID<5> , \pc_inc_two_ID<4> , \pc_inc_two_ID<3> ,
         \pc_inc_two_ID<2> , \pc_inc_two_ID<1> , \pc_inc_two_ID<0> , branch_id,
         haltID, jmp_r_ID, \rs<2> , \rs<1> , \rs<0> , \rd<2> , \rd<1> ,
         \rd<0> , \immID<15> , \immID<14> , \immID<13> , \immID<12> ,
         \immID<11> , \immID<10> , \immID<9> , \immID<8> , \immID<7> ,
         \immID<6> , \immID<5> , \immID<4> , \immID<3> , \immID<2> ,
         \immID<1> , \immID<0> , \displacementID<15> , \displacementID<14> ,
         \displacementID<13> , \displacementID<12> , \displacementID<11> ,
         \displacementID<10> , \displacementID<9> , \displacementID<8> ,
         \displacementID<7> , \displacementID<6> , \displacementID<5> ,
         \displacementID<4> , \displacementID<3> , \displacementID<2> ,
         \displacementID<1> , \displacementID<0> , \read1dataID<15> ,
         \read1dataID<14> , \read1dataID<13> , \read1dataID<12> ,
         \read1dataID<11> , \read1dataID<10> , \read1dataID<9> ,
         \read1dataID<8> , \read1dataID<7> , \read1dataID<6> ,
         \read1dataID<5> , \read1dataID<4> , \read1dataID<3> ,
         \read1dataID<2> , \read1dataID<1> , \read1dataID<0> ,
         \read2dataID<15> , \read2dataID<14> , \read2dataID<13> ,
         \read2dataID<12> , \read2dataID<11> , \read2dataID<10> ,
         \read2dataID<9> , \read2dataID<8> , \read2dataID<7> ,
         \read2dataID<6> , \read2dataID<5> , \read2dataID<4> ,
         \read2dataID<3> , \read2dataID<2> , \read2dataID<1> ,
         \read2dataID<0> , \r1_reg<2> , \r1_reg<1> , \r1_reg<0> , \r2_reg<2> ,
         \r2_reg<1> , \r2_reg<0> , \wb_r_wr<2> , \wb_r_wr<1> , \wb_r_wr<0> ,
         \regwritedata<15> , \regwritedata<14> , \regwritedata<13> ,
         \regwritedata<12> , \regwritedata<11> , \regwritedata<10> ,
         \regwritedata<9> , \regwritedata<8> , \regwritedata<7> ,
         \regwritedata<6> , \regwritedata<5> , \regwritedata<4> ,
         \regwritedata<3> , \regwritedata<2> , \regwritedata<1> ,
         \regwritedata<0> , regwrite, id_rs_v, id_rt_v, id_rd_v, \r_wr<2> ,
         \r_wr<1> , \r_wr<0> , fow_EXID_rs_ID, fow_MEMID_rs_ID, fow_EXID_rt_ID,
         fow_MEMID_rt_ID, \wr_aluOut<15> , \wr_aluOut<14> , \wr_aluOut<13> ,
         \wr_aluOut<12> , \wr_aluOut<11> , \wr_aluOut<10> , \wr_aluOut<9> ,
         \wr_aluOut<8> , \wr_aluOut<7> , \wr_aluOut<6> , \wr_aluOut<5> ,
         \wr_aluOut<4> , \wr_aluOut<3> , \wr_aluOut<2> , \wr_aluOut<1> ,
         \wr_aluOut<0> , \aluOut<15> , \aluOut<14> , \aluOut<13> ,
         \aluOut<12> , \aluOut<11> , \aluOut<10> , \aluOut<9> , \aluOut<8> ,
         \aluOut<7> , \aluOut<6> , \aluOut<5> , \aluOut<4> , \aluOut<3> ,
         \aluOut<2> , \aluOut<1> , \aluOut<0> , \rdEX<2> , \rdEX<1> ,
         \rdEX<0> , \rsEX<2> , \rsEX<1> , \rsEX<0> , \ex_r_wr<2> ,
         \ex_r_wr<1> , \ex_r_wr<0> , \read1dataEX<15> , \read1dataEX<14> ,
         \read1dataEX<13> , \read1dataEX<12> , \read1dataEX<11> ,
         \read1dataEX<10> , \read1dataEX<9> , \read1dataEX<8> ,
         \read1dataEX<7> , \read1dataEX<6> , \read1dataEX<5> ,
         \read1dataEX<4> , \read1dataEX<3> , \read1dataEX<2> ,
         \read1dataEX<1> , \read1dataEX<0> , \read2dataEX<15> ,
         \read2dataEX<14> , \read2dataEX<13> , \read2dataEX<12> ,
         \read2dataEX<11> , \read2dataEX<10> , \read2dataEX<9> ,
         \read2dataEX<8> , \read2dataEX<7> , \read2dataEX<6> ,
         \read2dataEX<5> , \read2dataEX<4> , \read2dataEX<3> ,
         \read2dataEX<2> , \read2dataEX<1> , \read2dataEX<0> , \immEX<15> ,
         \immEX<14> , \immEX<13> , \immEX<12> , \immEX<11> , \immEX<10> ,
         \immEX<9> , \immEX<8> , \immEX<7> , \immEX<6> , \immEX<5> ,
         \immEX<4> , \immEX<3> , \immEX<2> , \immEX<1> , \immEX<0> , ex_rd_v,
         haltEX, \pc_inc_two_EX<15> , \pc_inc_two_EX<14> , \pc_inc_two_EX<13> ,
         \pc_inc_two_EX<12> , \pc_inc_two_EX<11> , \pc_inc_two_EX<10> ,
         \pc_inc_two_EX<9> , \pc_inc_two_EX<8> , \pc_inc_two_EX<7> ,
         \pc_inc_two_EX<6> , \pc_inc_two_EX<5> , \pc_inc_two_EX<4> ,
         \pc_inc_two_EX<3> , \pc_inc_two_EX<2> , \pc_inc_two_EX<1> ,
         \pc_inc_two_EX<0> , fow_EXID_rs_EX, fow_MEMID_rs_EX, fow_EXID_rt_EX,
         fow_MEMID_rt_EX, \nx_pcEX<15> , \nx_pcEX<14> , \nx_pcEX<13> ,
         \nx_pcEX<12> , \nx_pcEX<11> , \nx_pcEX<10> , \nx_pcEX<9> ,
         \nx_pcEX<8> , \nx_pcEX<7> , \nx_pcEX<6> , \nx_pcEX<5> , \nx_pcEX<4> ,
         \nx_pcEX<3> , \nx_pcEX<2> , \nx_pcEX<1> , \nx_pcEX<0> ,
         \regwritedata_m<15> , \regwritedata_m<14> , \regwritedata_m<13> ,
         \regwritedata_m<12> , \regwritedata_m<11> , \regwritedata_m<10> ,
         \regwritedata_m<9> , \regwritedata_m<8> , \regwritedata_m<7> ,
         \regwritedata_m<6> , \regwritedata_m<5> , \regwritedata_m<4> ,
         \regwritedata_m<3> , \regwritedata_m<2> , \regwritedata_m<1> ,
         \regwritedata_m<0> , \forwarded_read2dataEX<15> ,
         \forwarded_read2dataEX<12> , \forwarded_read2dataEX<9> ,
         \forwarded_read2dataEX<8> , \forwarded_read2dataEX<5> ,
         \forwarded_read2dataEX<4> , alusrc, \opB<15> , \opB<13> , \opB<12> ,
         \opB<10> , \opB<2> , cin, \alu_op<2> , \alu_op<1> , \alu_op<0> , invA,
         invB, ofl, zero, N, P, c_out, \shamt<3> , \shamt<2> , \shamt<1> ,
         \shamt<0> , shift, slbi_EX, \rdMEM<2> , \rdMEM<1> , \rdMEM<0> ,
         \rsMEM<2> , \rsMEM<1> , \rsMEM<0> , \mem_r_wr<2> , \mem_r_wr<1> ,
         \mem_r_wr<0> , \instMEM_normal<15> , \instMEM_normal<14> ,
         \instMEM_normal<13> , \instMEM_normal<12> , \instMEM_normal<11> ,
         \instMEM_normal<10> , \instMEM_normal<9> , \instMEM_normal<8> ,
         \instMEM_normal<7> , \instMEM_normal<6> , \instMEM_normal<5> ,
         \instMEM_normal<4> , \instMEM_normal<3> , \instMEM_normal<2> ,
         \instMEM_normal<1> , \instMEM_normal<0> , \aluOutMEM<15> ,
         \aluOutMEM<14> , \aluOutMEM<13> , \aluOutMEM<12> , \aluOutMEM<11> ,
         \aluOutMEM<10> , \aluOutMEM<9> , \aluOutMEM<8> , \aluOutMEM<7> ,
         \aluOutMEM<6> , \aluOutMEM<5> , \aluOutMEM<4> , \aluOutMEM<3> ,
         \aluOutMEM<2> , \aluOutMEM<1> , \aluOutMEM<0> , \read1dataMEM<15> ,
         \read1dataMEM<14> , \read1dataMEM<13> , \read1dataMEM<12> ,
         \read1dataMEM<11> , \read1dataMEM<10> , \read1dataMEM<9> ,
         \read1dataMEM<8> , \read1dataMEM<7> , \read1dataMEM<6> ,
         \read1dataMEM<5> , \read1dataMEM<4> , \read1dataMEM<3> ,
         \read1dataMEM<2> , \read1dataMEM<1> , \read1dataMEM<0> ,
         \read2dataMEM<15> , \read2dataMEM<14> , \read2dataMEM<13> ,
         \read2dataMEM<12> , \read2dataMEM<11> , \read2dataMEM<10> ,
         \read2dataMEM<9> , \read2dataMEM<8> , \read2dataMEM<7> ,
         \read2dataMEM<6> , \read2dataMEM<5> , \read2dataMEM<4> ,
         \read2dataMEM<3> , \read2dataMEM<2> , \read2dataMEM<1> ,
         \read2dataMEM<0> , \immMEM<15> , \immMEM<14> , \immMEM<13> ,
         \immMEM<12> , \immMEM<11> , \immMEM<10> , \immMEM<9> , \immMEM<8> ,
         \immMEM<7> , \immMEM<6> , \immMEM<5> , \immMEM<4> , \immMEM<3> ,
         \immMEM<2> , \immMEM<1> , \immMEM<0> , \forwarded_read2dataMEM<15> ,
         \forwarded_read2dataMEM<14> , \forwarded_read2dataMEM<13> ,
         \forwarded_read2dataMEM<12> , \forwarded_read2dataMEM<11> ,
         \forwarded_read2dataMEM<10> , \forwarded_read2dataMEM<9> ,
         \forwarded_read2dataMEM<8> , \forwarded_read2dataMEM<7> ,
         \forwarded_read2dataMEM<6> , \forwarded_read2dataMEM<5> ,
         \forwarded_read2dataMEM<4> , \forwarded_read2dataMEM<3> ,
         \forwarded_read2dataMEM<2> , \forwarded_read2dataMEM<1> ,
         \forwarded_read2dataMEM<0> , \pc_inc_two_MEM<15> ,
         \pc_inc_two_MEM<14> , \pc_inc_two_MEM<13> , \pc_inc_two_MEM<12> ,
         \pc_inc_two_MEM<11> , \pc_inc_two_MEM<10> , \pc_inc_two_MEM<9> ,
         \pc_inc_two_MEM<8> , \pc_inc_two_MEM<7> , \pc_inc_two_MEM<6> ,
         \pc_inc_two_MEM<5> , \pc_inc_two_MEM<4> , \pc_inc_two_MEM<3> ,
         \pc_inc_two_MEM<2> , \pc_inc_two_MEM<1> , \pc_inc_two_MEM<0> , oflMEM,
         c_outMEM, zeroMEM, NMEM, PMEM, mem_rd_v, slbi_MEM, \nx_pcMEM<15> ,
         \nx_pcMEM<14> , \nx_pcMEM<13> , \nx_pcMEM<12> , \nx_pcMEM<11> ,
         \nx_pcMEM<10> , \nx_pcMEM<9> , \nx_pcMEM<8> , \nx_pcMEM<7> ,
         \nx_pcMEM<6> , \nx_pcMEM<5> , \nx_pcMEM<4> , \nx_pcMEM<3> ,
         \nx_pcMEM<2> , \nx_pcMEM<1> , \nx_pcMEM<0> , memread, memwrite,
         memtoreg_m, ld_imm_m, compareS_m, btr_m, regdst_m, \mem_out<15> ,
         \mem_out<14> , \mem_out<13> , \mem_out<12> , \mem_out<11> ,
         \mem_out<10> , \mem_out<9> , \mem_out<8> , \mem_out<7> , \mem_out<6> ,
         \mem_out<5> , \mem_out<4> , \mem_out<3> , \mem_out<2> , \mem_out<1> ,
         \mem_out<0> , memDone, memStall, \rdWB<2> , \rdWB<1> , \rdWB<0> ,
         \rsWB<2> , \rsWB<1> , \rsWB<0> , \instWB_normal<15> ,
         \instWB_normal<14> , \instWB_normal<13> , \instWB_normal<12> ,
         \instWB_normal<11> , \instWB_normal<10> , \instWB_normal<9> ,
         \instWB_normal<8> , \instWB_normal<7> , \instWB_normal<6> ,
         \instWB_normal<5> , \instWB_normal<4> , \instWB_normal<3> ,
         \instWB_normal<2> , \instWB_normal<1> , \instWB_normal<0> ,
         \aluOutWB<15> , \aluOutWB<14> , \aluOutWB<13> , \aluOutWB<12> ,
         \aluOutWB<11> , \aluOutWB<10> , \aluOutWB<9> , \aluOutWB<8> ,
         \aluOutWB<7> , \aluOutWB<6> , \aluOutWB<5> , \aluOutWB<4> ,
         \aluOutWB<3> , \aluOutWB<2> , \aluOutWB<1> , \aluOutWB<0> ,
         \mem_outWB<15> , \mem_outWB<14> , \mem_outWB<13> , \mem_outWB<12> ,
         \mem_outWB<11> , \mem_outWB<10> , \mem_outWB<9> , \mem_outWB<8> ,
         \mem_outWB<7> , \mem_outWB<6> , \mem_outWB<5> , \mem_outWB<4> ,
         \mem_outWB<3> , \mem_outWB<2> , \mem_outWB<1> , \mem_outWB<0> ,
         \immWB<15> , \immWB<14> , \immWB<13> , \immWB<12> , \immWB<11> ,
         \immWB<10> , \immWB<9> , \immWB<8> , \immWB<7> , \immWB<6> ,
         \immWB<5> , \immWB<4> , \immWB<3> , \immWB<2> , \immWB<1> ,
         \immWB<0> , \pc_inc_two_WB<15> , \pc_inc_two_WB<14> ,
         \pc_inc_two_WB<13> , \pc_inc_two_WB<12> , \pc_inc_two_WB<11> ,
         \pc_inc_two_WB<10> , \pc_inc_two_WB<9> , \pc_inc_two_WB<8> ,
         \pc_inc_two_WB<7> , \pc_inc_two_WB<6> , \pc_inc_two_WB<5> ,
         \pc_inc_two_WB<4> , \pc_inc_two_WB<3> , \pc_inc_two_WB<2> ,
         \pc_inc_two_WB<1> , \pc_inc_two_WB<0> , oflWB, zeroWB, NWB, PWB,
         c_outWB, slbi_WB, memtoreg, ld_imm, compareS, btr, writeR7, regdst,
         n8, n9, n65, n69, n71, n73, n75, n77, n79, n81, n83, n85, n87, n89,
         n91, n96, n98, n124, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207;

  dff_665 stal ( .q(), .d(stall), .clk(clk), .rst(n986) );
  reg1_26 instMemDoneReg ( .d(n746), .q(instMemDone_q), .clk(clk), .rst(n985), 
        .en(1'b1) );
  reg16_36 instIFReg ( .read({\instIF_q<15> , \instIF_q<14> , \instIF_q<13> , 
        \instIF_q<12> , \instIF_q<11> , \instIF_q<10> , \instIF_q<9> , 
        \instIF_q<8> , \instIF_q<7> , \instIF_q<6> , \instIF_q<5> , 
        \instIF_q<4> , \instIF_q<3> , \instIF_q<2> , \instIF_q<1> , 
        \instIF_q<0> }), .write({n9, n8, n828, n826, n675, n824, n822, n820, 
        n818, n816, n814, n812, n810, n808, n806, n804}), .wr_en(n1204), .rst(
        n985), .clk(clk) );
  IF_control ifcont ( .Jump(jump_IF), .Branch(branch_if), .jmp_r(), .opcode({
        n9, n8, n828, n826, n675}) );
  pc prog_c ( .branch_if(branch_if), .pc_inc_two({\pc_inc_two<15> , 
        \pc_inc_two<14> , \pc_inc_two<13> , \pc_inc_two<12> , \pc_inc_two<11> , 
        \pc_inc_two<10> , \pc_inc_two<9> , \pc_inc_two<8> , \pc_inc_two<7> , 
        \pc_inc_two<6> , \pc_inc_two<5> , \pc_inc_two<4> , \pc_inc_two<3> , 
        \pc_inc_two<2> , \pc_inc_two<1> , \pc_inc_two<0> }), .jmp_r(1'b0), 
        .en(pc_en), .clk(clk), .rst(n986), .jump(jump_EX), .inst({n9, n8, n828, 
        n826, n675, n824, n822, n820, n818, n816, n814, n812, n810, n808, n806, 
        n804}), .addr({\addr<15> , \addr<14> , \addr<13> , \addr<12> , 
        \addr<11> , \addr<10> , \addr<9> , \addr<8> , \addr<7> , \addr<6> , 
        \addr<5> , \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), 
        .branch(branch_ex), .rs({\forwarded_read1dataEX<15> , n946, 
        \forwarded_read1dataEX<13> , \forwarded_read1dataEX<12> , n277, n243, 
        \forwarded_read1dataEX<9> , n926, n908, n637, 
        \forwarded_read1dataEX<5> , n640, n633, n544, n962, n240}), .pc_nx({
        \pc_nx<15> , \pc_nx<14> , \pc_nx<13> , \pc_nx<12> , \pc_nx<11> , 
        \pc_nx<10> , \pc_nx<9> , \pc_nx<8> , \pc_nx<7> , \pc_nx<6> , 
        \pc_nx<5> , \pc_nx<4> , \pc_nx<3> , \pc_nx<2> , \pc_nx<1> , \pc_nx<0> }), .EX_inst({n194, n218, n181, n198, n226, \instEX_normal<10> , 
        \instEX_normal<9> , \instEX_normal<8> , \instEX_normal<7> , 
        \instEX_normal<6> , \instEX_normal<5> , \instEX_normal<4> , 
        \instEX_normal<3> , \instEX_normal<2> , \instEX_normal<1> , 
        \instEX_normal<0> }), .br_ctl(br_ctl) );
  mem_system inst_mem ( .DataOut({\instIF_normal<15> , \instIF_normal<14> , 
        \instIF_normal<13> , \instIF_normal<12> , \instIF_normal<11> , 
        \instIF_normal<10> , \instIF_normal<9> , \instIF_normal<8> , 
        \instIF_normal<7> , \instIF_normal<6> , \instIF_normal<5> , 
        \instIF_normal<4> , \instIF_normal<3> , \instIF_normal<2> , 
        \instIF_normal<1> , \instIF_normal<0> }), .Done(instMemDone), .Stall(
        instMemStall), .CacheHit(), .err(IcacheErr), .Addr({\addr<15> , 
        \addr<14> , \addr<13> , \addr<12> , \addr<11> , \addr<10> , \addr<9> , 
        \addr<8> , \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , 
        \addr<2> , \addr<1> , \addr<0> }), .DataIn({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Rd(_3_net_), .Wr(1'b0), .clk(clk), .rst(rst) );
  reg16_init IFID ( .read({\instID<15> , \instID<14> , \instID<13> , 
        \instID<12> , \instID<11> , \instID<10> , \instID<9> , \instID<8> , 
        \instID<7> , \instID<6> , \instID<5> , \instID<4> , \instID<3> , 
        \instID<2> , \instID<1> , \instID<0> }), .write({\wr_instIF<15> , 
        \wr_instIF<14> , \wr_instIF<13> , \wr_instIF<12> , \wr_instIF<11> , 
        \wr_instIF<10> , \wr_instIF<9> , \wr_instIF<8> , \wr_instIF<7> , 
        \wr_instIF<6> , \wr_instIF<5> , \wr_instIF<4> , \wr_instIF<3> , 
        \wr_instIF<2> , \wr_instIF<1> , \wr_instIF<0> }), .wr_en(n988), .rst(
        n914), .clk(clk) );
  reg16_35 nx_pcid ( .read({\nx_pcID<15> , \nx_pcID<14> , \nx_pcID<13> , 
        \nx_pcID<12> , \nx_pcID<11> , \nx_pcID<10> , \nx_pcID<9> , 
        \nx_pcID<8> , \nx_pcID<7> , \nx_pcID<6> , \nx_pcID<5> , \nx_pcID<4> , 
        \nx_pcID<3> , \nx_pcID<2> , \nx_pcID<1> , \nx_pcID<0> }), .write({
        \pc_nx<15> , \pc_nx<14> , \pc_nx<13> , \pc_nx<12> , \pc_nx<11> , 
        \pc_nx<10> , \pc_nx<9> , \pc_nx<8> , \pc_nx<7> , \pc_nx<6> , 
        \pc_nx<5> , \pc_nx<4> , \pc_nx<3> , \pc_nx<2> , \pc_nx<1> , \pc_nx<0> }), .wr_en(n1007), .rst(n985), .clk(clk) );
  reg16_34 pc_inc_twoid ( .read({\pc_inc_two_ID<15> , \pc_inc_two_ID<14> , 
        \pc_inc_two_ID<13> , \pc_inc_two_ID<12> , \pc_inc_two_ID<11> , 
        \pc_inc_two_ID<10> , \pc_inc_two_ID<9> , \pc_inc_two_ID<8> , 
        \pc_inc_two_ID<7> , \pc_inc_two_ID<6> , \pc_inc_two_ID<5> , 
        \pc_inc_two_ID<4> , \pc_inc_two_ID<3> , \pc_inc_two_ID<2> , 
        \pc_inc_two_ID<1> , \pc_inc_two_ID<0> }), .write({\pc_inc_two<15> , 
        \pc_inc_two<14> , \pc_inc_two<13> , \pc_inc_two<12> , \pc_inc_two<11> , 
        \pc_inc_two<10> , \pc_inc_two<9> , \pc_inc_two<8> , \pc_inc_two<7> , 
        \pc_inc_two<6> , \pc_inc_two<5> , \pc_inc_two<4> , \pc_inc_two<3> , 
        \pc_inc_two<2> , \pc_inc_two<1> , \pc_inc_two<0> }), .wr_en(n988), 
        .rst(n986), .clk(clk) );
  reg1_25 branchid ( .d(n518), .q(branch_id), .clk(clk), .rst(n986), .en(n988)
         );
  reg1_24 jumpid ( .d(n516), .q(jump_ID), .clk(clk), .rst(n986), .en(n988) );
  ID_control idcont ( .Rt_Rd(), .Halt(haltID), .jmp_r(jmp_r_ID), .opcode({
        \instID<15> , \instID<14> , \instID<13> , \instID<12> , \instID<11> })
         );
  decoder inst_decode ( .inst({\instID<15> , \instID<14> , \instID<13> , 
        \instID<12> , \instID<11> , \instID<10> , \instID<9> , \instID<8> , 
        \instID<7> , \instID<6> , \instID<5> , \instID<4> , \instID<3> , 
        \instID<2> , \instID<1> , \instID<0> }), .rt(), .rs({\rs<2> , \rs<1> , 
        \rs<0> }), .rd({\rd<2> , \rd<1> , \rd<0> }), .imm({\immID<15> , 
        \immID<14> , \immID<13> , \immID<12> , \immID<11> , \immID<10> , 
        \immID<9> , \immID<8> , \immID<7> , \immID<6> , \immID<5> , \immID<4> , 
        \immID<3> , \immID<2> , \immID<1> , \immID<0> }), .displacement({
        \displacementID<15> , \displacementID<14> , \displacementID<13> , 
        \displacementID<12> , \displacementID<11> , \displacementID<10> , 
        \displacementID<9> , \displacementID<8> , \displacementID<7> , 
        \displacementID<6> , \displacementID<5> , \displacementID<4> , 
        \displacementID<3> , \displacementID<2> , \displacementID<1> , 
        \displacementID<0> }) );
  rf_bypass regfile ( .read1data({\read1dataID<15> , \read1dataID<14> , 
        \read1dataID<13> , \read1dataID<12> , \read1dataID<11> , 
        \read1dataID<10> , \read1dataID<9> , \read1dataID<8> , 
        \read1dataID<7> , \read1dataID<6> , \read1dataID<5> , \read1dataID<4> , 
        \read1dataID<3> , \read1dataID<2> , \read1dataID<1> , \read1dataID<0> }), .read2data({\read2dataID<15> , \read2dataID<14> , \read2dataID<13> , 
        \read2dataID<12> , \read2dataID<11> , \read2dataID<10> , 
        \read2dataID<9> , \read2dataID<8> , \read2dataID<7> , \read2dataID<6> , 
        \read2dataID<5> , \read2dataID<4> , \read2dataID<3> , \read2dataID<2> , 
        \read2dataID<1> , \read2dataID<0> }), .err(rf_bypass_err), .clk(clk), 
        .rst(n985), .read1regsel({\r1_reg<2> , \r1_reg<1> , \r1_reg<0> }), 
        .read2regsel({\r2_reg<2> , \r2_reg<1> , \r2_reg<0> }), .writeregsel({
        \wb_r_wr<2> , \wb_r_wr<1> , \wb_r_wr<0> }), .writedata({n960, n974, 
        n217, n937, n909, n964, n966, n212, n197, n931, n973, n983, n972, n231, 
        n204, n982}), .write(regwrite) );
  reg_control regctl ( .rs_v(id_rs_v), .rt_v(id_rt_v), .rd_v(id_rd_v), 
        .r1_reg({\r1_reg<2> , \r1_reg<1> , \r1_reg<0> }), .r2_reg({\r2_reg<2> , 
        \r2_reg<1> , \r2_reg<0> }), .r_wr({\r_wr<2> , \r_wr<1> , \r_wr<0> }), 
        .inst({\instID<15> , \instID<14> , \instID<13> , \instID<12> , 
        \instID<11> , \instID<10> , \instID<9> , \instID<8> , \instID<7> , 
        \instID<6> , \instID<5> , \instID<4> , \instID<3> , \instID<2> , 
        \instID<1> , \instID<0> }) );
  reg3_8 rdex ( .read({\rdEX<2> , \rdEX<1> , \rdEX<0> }), .write({n514, n512, 
        n510}), .wr_en(n1007), .rst(n985), .clk(clk) );
  reg3_7 rsex ( .read({\rsEX<2> , \rsEX<1> , \rsEX<0> }), .write({n508, n506, 
        n504}), .wr_en(n989), .rst(n985), .clk(clk) );
  reg3_6 rwrex ( .read({\ex_r_wr<2> , \ex_r_wr<1> , \ex_r_wr<0> }), .write({
        n502, n500, n498}), .wr_en(n988), .rst(n986), .clk(clk) );
  reg16_33 instex ( .read({\instEX_normal<15> , \instEX_normal<14> , 
        \instEX_normal<13> , \instEX_normal<12> , \instEX_normal<11> , 
        \instEX_normal<10> , \instEX_normal<9> , \instEX_normal<8> , 
        \instEX_normal<7> , \instEX_normal<6> , \instEX_normal<5> , 
        \instEX_normal<4> , \instEX_normal<3> , \instEX_normal<2> , 
        \instEX_normal<1> , \instEX_normal<0> }), .write({n496, n494, n492, 
        n273, n681, n490, n488, n486, n484, n482, n480, n478, n476, n474, n472, 
        n470}), .wr_en(n988), .rst(n986), .clk(clk) );
  reg16_32 read1dataex ( .read({\read1dataEX<15> , \read1dataEX<14> , 
        \read1dataEX<13> , \read1dataEX<12> , \read1dataEX<11> , 
        \read1dataEX<10> , \read1dataEX<9> , \read1dataEX<8> , 
        \read1dataEX<7> , \read1dataEX<6> , \read1dataEX<5> , \read1dataEX<4> , 
        \read1dataEX<3> , \read1dataEX<2> , \read1dataEX<1> , \read1dataEX<0> }), .write({n468, n466, n464, n462, n460, n458, n456, n454, n452, n450, n448, 
        n446, n444, n442, n440, n438}), .wr_en(n1007), .rst(n985), .clk(clk)
         );
  reg16_31 read2dataex ( .read({\read2dataEX<15> , \read2dataEX<14> , 
        \read2dataEX<13> , \read2dataEX<12> , \read2dataEX<11> , 
        \read2dataEX<10> , \read2dataEX<9> , \read2dataEX<8> , 
        \read2dataEX<7> , \read2dataEX<6> , \read2dataEX<5> , \read2dataEX<4> , 
        \read2dataEX<3> , \read2dataEX<2> , \read2dataEX<1> , \read2dataEX<0> }), .write({n436, n434, n432, n430, n428, n426, n424, n422, n420, n418, n416, 
        n414, n412, n410, n408, n406}), .wr_en(n1007), .rst(n986), .clk(clk)
         );
  reg16_30 immex ( .read({\immEX<15> , \immEX<14> , \immEX<13> , \immEX<12> , 
        \immEX<11> , \immEX<10> , \immEX<9> , \immEX<8> , \immEX<7> , 
        \immEX<6> , \immEX<5> , \immEX<4> , \immEX<3> , \immEX<2> , \immEX<1> , 
        \immEX<0> }), .write({n669, n403, n669, n403, n403, n669, n669, n403, 
        n402, n400, n398, n396, n394, n392, n390, n388}), .wr_en(n1007), .rst(
        n985), .clk(clk) );
  reg16_29 disex ( .read(), .write({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n386, n384, 
        n382, n380, n378, n376, n374, n372, n370, n368, n366}), .wr_en(n988), 
        .rst(n986), .clk(clk) );
  reg1_23 rdexv ( .d(n364), .q(ex_rd_v), .clk(clk), .rst(n986), .en(n1007) );
  reg1_22 haltex ( .d(n362), .q(haltEX), .clk(clk), .rst(n985), .en(n1007) );
  reg16_28 pc_inc_twoex ( .read({\pc_inc_two_EX<15> , \pc_inc_two_EX<14> , 
        \pc_inc_two_EX<13> , \pc_inc_two_EX<12> , \pc_inc_two_EX<11> , 
        \pc_inc_two_EX<10> , \pc_inc_two_EX<9> , \pc_inc_two_EX<8> , 
        \pc_inc_two_EX<7> , \pc_inc_two_EX<6> , \pc_inc_two_EX<5> , 
        \pc_inc_two_EX<4> , \pc_inc_two_EX<3> , \pc_inc_two_EX<2> , 
        \pc_inc_two_EX<1> , \pc_inc_two_EX<0> }), .write({n360, n358, n356, 
        n354, n352, n350, n348, n346, n344, n342, n340, n338, n336, n271, n334, 
        n269}), .wr_en(n989), .rst(n985), .clk(clk) );
  reg1_21 ex_rs ( .d(n267), .q(fow_EXID_rs_EX), .clk(clk), .rst(n986), .en(
        n989) );
  reg1_20 mem_rs ( .d(n332), .q(fow_MEMID_rs_EX), .clk(clk), .rst(n985), .en(
        n988) );
  reg1_19 ex_rt ( .d(n330), .q(fow_EXID_rt_EX), .clk(clk), .rst(n986), .en(
        n988) );
  reg1_18 mem_rt ( .d(n265), .q(fow_MEMID_rt_EX), .clk(clk), .rst(n985), .en(
        n1007) );
  reg1_17 jmp_rex ( .d(n328), .q(), .clk(clk), .rst(n986), .en(n1007) );
  reg16_27 nx_pcex ( .read({\nx_pcEX<15> , \nx_pcEX<14> , \nx_pcEX<13> , 
        \nx_pcEX<12> , \nx_pcEX<11> , \nx_pcEX<10> , \nx_pcEX<9> , 
        \nx_pcEX<8> , \nx_pcEX<7> , \nx_pcEX<6> , \nx_pcEX<5> , \nx_pcEX<4> , 
        \nx_pcEX<3> , \nx_pcEX<2> , \nx_pcEX<1> , \nx_pcEX<0> }), .write({n326, 
        n263, n324, n261, n322, n259, n320, n257, n318, n255, n316, n253, n314, 
        n251, n312, n249}), .wr_en(n989), .rst(n986), .clk(clk) );
  reg16_26 aluO_ex ( .read(), .write({\wr_aluOut<15> , \wr_aluOut<14> , 
        \wr_aluOut<13> , \wr_aluOut<12> , \wr_aluOut<11> , \wr_aluOut<10> , 
        \wr_aluOut<9> , \wr_aluOut<8> , \wr_aluOut<7> , \wr_aluOut<6> , 
        \wr_aluOut<5> , \wr_aluOut<4> , \wr_aluOut<3> , \wr_aluOut<2> , 
        \wr_aluOut<1> , \wr_aluOut<0> }), .wr_en(n1007), .rst(n985), .clk(clk)
         );
  reg1_16 branchex ( .d(n247), .q(branch_ex), .clk(clk), .rst(n985), .en(n989)
         );
  reg1_15 jumpex ( .d(n245), .q(jump_EX), .clk(clk), .rst(n986), .en(n989) );
  EX_control excont ( .ALUOp(), .ALUSrc(alusrc), .wr_r7(), .compareS_EX(), 
        .opcode({\instEX_normal<15> , \instEX_normal<14> , \instEX_normal<13> , 
        n236, n226}) );
  alu ALU ( .A({n882, n206, n223, \forwarded_read1dataEX<12> , n211, n243, 
        n902, \forwarded_read1dataEX<8> , n188, n636, 
        \forwarded_read1dataEX<5> , n639, n633, n868, n303, n668}), .B({
        \opB<15> , n873, \opB<13> , \opB<12> , n216, \opB<10> , n295, n872, 
        n238, n630, n242, n870, n213, \opB<2> , n1207, n228}), .Cin(cin), .Op(
        {\alu_op<2> , \alu_op<1> , \alu_op<0> }), .invA(invA), .invB(invB), 
        .sign(1'b1), .Out({\aluOut<15> , \aluOut<14> , \aluOut<13> , 
        \aluOut<12> , \aluOut<11> , \aluOut<10> , \aluOut<9> , \aluOut<8> , 
        \aluOut<7> , \aluOut<6> , \aluOut<5> , \aluOut<4> , \aluOut<3> , 
        \aluOut<2> , \aluOut<1> , \aluOut<0> }), .Ofl(ofl), .Z(zero), .N(N), 
        .P(P), .c_out(c_out) );
  alu_control a_c ( .alu_op({\alu_op<2> , \alu_op<1> , \alu_op<0> }), .inv_a(
        invA), .inv_b(invB), .cin(cin), .shamt({\shamt<3> , \shamt<2> , 
        \shamt<1> , \shamt<0> }), .flip_1(), .flip_2(), .shift(shift), .SLBI(
        slbi_EX), .opcode({\instEX_normal<15> , \instEX_normal<14> , 
        \instEX_normal<13> , \instEX_normal<12> , \instEX_normal<11> }), 
        .func({\instEX_normal<1> , \instEX_normal<0> }), .immd({
        \instEX_normal<3> , \instEX_normal<2> , \instEX_normal<1> , 
        \instEX_normal<0> }) );
  reg3_5 rdmem ( .read({\rdMEM<2> , \rdMEM<1> , \rdMEM<0> }), .write({
        \rdEX<2> , \rdEX<1> , \rdEX<0> }), .wr_en(n988), .rst(n986), .clk(clk)
         );
  reg3_4 rsmem ( .read({\rsMEM<2> , \rsMEM<1> , \rsMEM<0> }), .write({
        \rsEX<2> , \rsEX<1> , \rsEX<0> }), .wr_en(n1007), .rst(n986), .clk(clk) );
  reg3_3 rwrmem ( .read({\mem_r_wr<2> , \mem_r_wr<1> , \mem_r_wr<0> }), 
        .write({\ex_r_wr<2> , \ex_r_wr<1> , \ex_r_wr<0> }), .wr_en(n1007), 
        .rst(n986), .clk(clk) );
  reg16_25 instM ( .read({\instMEM_normal<15> , \instMEM_normal<14> , 
        \instMEM_normal<13> , \instMEM_normal<12> , \instMEM_normal<11> , 
        \instMEM_normal<10> , \instMEM_normal<9> , \instMEM_normal<8> , 
        \instMEM_normal<7> , \instMEM_normal<6> , \instMEM_normal<5> , 
        \instMEM_normal<4> , \instMEM_normal<3> , \instMEM_normal<2> , 
        \instMEM_normal<1> , \instMEM_normal<0> }), .write({n194, n218, n181, 
        n198, n226, \instEX_normal<10> , \instEX_normal<9> , 
        \instEX_normal<8> , \instEX_normal<7> , \instEX_normal<6> , 
        \instEX_normal<5> , \instEX_normal<4> , \instEX_normal<3> , 
        \instEX_normal<2> , \instEX_normal<1> , \instEX_normal<0> }), .wr_en(
        n988), .rst(n986), .clk(clk) );
  reg16_24 aluOutM ( .read({\aluOutMEM<15> , \aluOutMEM<14> , \aluOutMEM<13> , 
        \aluOutMEM<12> , \aluOutMEM<11> , \aluOutMEM<10> , \aluOutMEM<9> , 
        \aluOutMEM<8> , \aluOutMEM<7> , \aluOutMEM<6> , \aluOutMEM<5> , 
        \aluOutMEM<4> , \aluOutMEM<3> , \aluOutMEM<2> , \aluOutMEM<1> , 
        \aluOutMEM<0> }), .write({\aluOut<15> , \aluOut<14> , n938, n920, n956, 
        n933, n916, \aluOut<8> , \aluOut<7> , \aluOut<6> , n935, n897, 
        \aluOut<3> , \aluOut<2> , n894, \aluOut<0> }), .wr_en(n988), .rst(n986), .clk(clk) );
  reg16_23 read1dataM ( .read({\read1dataMEM<15> , \read1dataMEM<14> , 
        \read1dataMEM<13> , \read1dataMEM<12> , \read1dataMEM<11> , 
        \read1dataMEM<10> , \read1dataMEM<9> , \read1dataMEM<8> , 
        \read1dataMEM<7> , \read1dataMEM<6> , \read1dataMEM<5> , 
        \read1dataMEM<4> , \read1dataMEM<3> , \read1dataMEM<2> , 
        \read1dataMEM<1> , \read1dataMEM<0> }), .write({
        \forwarded_read1dataEX<15> , n947, n853, \forwarded_read1dataEX<12> , 
        n277, n243, n755, n200, n879, n874, \forwarded_read1dataEX<5> , n639, 
        n876, n871, n903, n761}), .wr_en(n988), .rst(n986), .clk(clk) );
  reg16_22 read2dataM ( .read({\read2dataMEM<15> , \read2dataMEM<14> , 
        \read2dataMEM<13> , \read2dataMEM<12> , \read2dataMEM<11> , 
        \read2dataMEM<10> , \read2dataMEM<9> , \read2dataMEM<8> , 
        \read2dataMEM<7> , \read2dataMEM<6> , \read2dataMEM<5> , 
        \read2dataMEM<4> , \read2dataMEM<3> , \read2dataMEM<2> , 
        \read2dataMEM<1> , \read2dataMEM<0> }), .write({\opB<15> , n873, n854, 
        \opB<12> , n284, \opB<10> , n185, n872, n672, n631, n763, n950, n910, 
        n205, n783, n875}), .wr_en(n988), .rst(n986), .clk(clk) );
  reg16_21 immM ( .read({\immMEM<15> , \immMEM<14> , \immMEM<13> , 
        \immMEM<12> , \immMEM<11> , \immMEM<10> , \immMEM<9> , \immMEM<8> , 
        \immMEM<7> , \immMEM<6> , \immMEM<5> , \immMEM<4> , \immMEM<3> , 
        \immMEM<2> , \immMEM<1> , \immMEM<0> }), .write({\immEX<15> , 
        \immEX<14> , \immEX<13> , \immEX<12> , \immEX<11> , \immEX<10> , 
        \immEX<9> , \immEX<8> , \immEX<7> , \immEX<6> , \immEX<5> , \immEX<4> , 
        \immEX<3> , \immEX<2> , \immEX<1> , \immEX<0> }), .wr_en(n989), .rst(
        n986), .clk(clk) );
  reg16_20 reg_forwarded_read2dataMEM ( .read({\forwarded_read2dataMEM<15> , 
        \forwarded_read2dataMEM<14> , \forwarded_read2dataMEM<13> , 
        \forwarded_read2dataMEM<12> , \forwarded_read2dataMEM<11> , 
        \forwarded_read2dataMEM<10> , \forwarded_read2dataMEM<9> , 
        \forwarded_read2dataMEM<8> , \forwarded_read2dataMEM<7> , 
        \forwarded_read2dataMEM<6> , \forwarded_read2dataMEM<5> , 
        \forwarded_read2dataMEM<4> , \forwarded_read2dataMEM<3> , 
        \forwarded_read2dataMEM<2> , \forwarded_read2dataMEM<1> , 
        \forwarded_read2dataMEM<0> }), .write({\forwarded_read2dataEX<15> , 
        n765, n767, \forwarded_read2dataEX<12> , n769, n771, n756, 
        \forwarded_read2dataEX<8> , n773, n757, n758, n759, n775, n777, n779, 
        n781}), .wr_en(n988), .rst(n986), .clk(clk) );
  reg16_19 pc_inc_twomem ( .read({\pc_inc_two_MEM<15> , \pc_inc_two_MEM<14> , 
        \pc_inc_two_MEM<13> , \pc_inc_two_MEM<12> , \pc_inc_two_MEM<11> , 
        \pc_inc_two_MEM<10> , \pc_inc_two_MEM<9> , \pc_inc_two_MEM<8> , 
        \pc_inc_two_MEM<7> , \pc_inc_two_MEM<6> , \pc_inc_two_MEM<5> , 
        \pc_inc_two_MEM<4> , \pc_inc_two_MEM<3> , \pc_inc_two_MEM<2> , 
        \pc_inc_two_MEM<1> , \pc_inc_two_MEM<0> }), .write({
        \pc_inc_two_EX<15> , \pc_inc_two_EX<14> , \pc_inc_two_EX<13> , 
        \pc_inc_two_EX<12> , \pc_inc_two_EX<11> , \pc_inc_two_EX<10> , 
        \pc_inc_two_EX<9> , \pc_inc_two_EX<8> , \pc_inc_two_EX<7> , 
        \pc_inc_two_EX<6> , \pc_inc_two_EX<5> , \pc_inc_two_EX<4> , 
        \pc_inc_two_EX<3> , \pc_inc_two_EX<2> , \pc_inc_two_EX<1> , 
        \pc_inc_two_EX<0> }), .wr_en(n989), .rst(n985), .clk(clk) );
  reg1_14 oflM ( .d(ofl), .q(oflMEM), .clk(clk), .rst(n985), .en(n988) );
  reg1_13 c_outM ( .d(c_out), .q(c_outMEM), .clk(clk), .rst(n986), .en(n1007)
         );
  reg1_12 zeroM ( .d(zero), .q(zeroMEM), .clk(clk), .rst(n985), .en(n989) );
  reg1_11 NM ( .d(N), .q(NMEM), .clk(clk), .rst(n986), .en(n989) );
  reg1_10 PM ( .d(P), .q(PMEM), .clk(clk), .rst(n985), .en(n1007) );
  reg1_9 rdmemv ( .d(ex_rd_v), .q(mem_rd_v), .clk(clk), .rst(n985), .en(n989)
         );
  reg1_8 haltmem ( .d(haltEX), .q(haltMEM), .clk(clk), .rst(n985), .en(n1007)
         );
  reg1_7 slbimem ( .d(slbi_EX), .q(slbi_MEM), .clk(clk), .rst(n985), .en(n988)
         );
  reg16_18 nx_pcmem ( .read({\nx_pcMEM<15> , \nx_pcMEM<14> , \nx_pcMEM<13> , 
        \nx_pcMEM<12> , \nx_pcMEM<11> , \nx_pcMEM<10> , \nx_pcMEM<9> , 
        \nx_pcMEM<8> , \nx_pcMEM<7> , \nx_pcMEM<6> , \nx_pcMEM<5> , 
        \nx_pcMEM<4> , \nx_pcMEM<3> , \nx_pcMEM<2> , \nx_pcMEM<1> , 
        \nx_pcMEM<0> }), .write({\nx_pcEX<15> , \nx_pcEX<14> , \nx_pcEX<13> , 
        \nx_pcEX<12> , \nx_pcEX<11> , \nx_pcEX<10> , \nx_pcEX<9> , 
        \nx_pcEX<8> , \nx_pcEX<7> , \nx_pcEX<6> , \nx_pcEX<5> , \nx_pcEX<4> , 
        \nx_pcEX<3> , \nx_pcEX<2> , \nx_pcEX<1> , \nx_pcEX<0> }), .wr_en(n989), 
        .rst(n986), .clk(clk) );
  MEM_control memcont ( .MemRead(memread), .MemWrite(memwrite), .opcode({n952, 
        n917, n928, n957, n941}) );
  WB_control_1 mem_wbcntl ( .MemtoReg(memtoreg_m), .RegWrite(), .ld_imm(
        ld_imm_m), .compareS(compareS_m), .btr(btr_m), .writeR7(), .RegDst(
        regdst_m), .opcode({\instMEM_normal<15> , \instMEM_normal<14> , 
        \instMEM_normal<13> , \instMEM_normal<12> , \instMEM_normal<11> }) );
  mem_system d_mem ( .DataOut({\mem_out<15> , \mem_out<14> , \mem_out<13> , 
        \mem_out<12> , \mem_out<11> , \mem_out<10> , \mem_out<9> , 
        \mem_out<8> , \mem_out<7> , \mem_out<6> , \mem_out<5> , \mem_out<4> , 
        \mem_out<3> , \mem_out<2> , \mem_out<1> , \mem_out<0> }), .Done(
        memDone), .Stall(memStall), .CacheHit(), .err(DcacheErr), .Addr({
        \aluOutMEM<15> , \aluOutMEM<14> , \aluOutMEM<13> , \aluOutMEM<12> , 
        \aluOutMEM<11> , \aluOutMEM<10> , \aluOutMEM<9> , \aluOutMEM<8> , 
        \aluOutMEM<7> , \aluOutMEM<6> , \aluOutMEM<5> , \aluOutMEM<4> , 
        \aluOutMEM<3> , \aluOutMEM<2> , \aluOutMEM<1> , \aluOutMEM<0> }), 
        .DataIn({\forwarded_read2dataMEM<15> , \forwarded_read2dataMEM<14> , 
        \forwarded_read2dataMEM<13> , \forwarded_read2dataMEM<12> , 
        \forwarded_read2dataMEM<11> , \forwarded_read2dataMEM<10> , 
        \forwarded_read2dataMEM<9> , \forwarded_read2dataMEM<8> , 
        \forwarded_read2dataMEM<7> , \forwarded_read2dataMEM<6> , 
        \forwarded_read2dataMEM<5> , \forwarded_read2dataMEM<4> , 
        \forwarded_read2dataMEM<3> , \forwarded_read2dataMEM<2> , 
        \forwarded_read2dataMEM<1> , \forwarded_read2dataMEM<0> }), .Rd(
        memread), .Wr(memwrite), .clk(clk), .rst(rst) );
  mf_data mdata ( .rd({\rdMEM<2> , \rdMEM<1> , \rdMEM<0> }), .rs({\rsMEM<2> , 
        \rsMEM<1> , \rsMEM<0> }), .regdst(regdst_m), .memtoreg(memtoreg_m), 
        .slbi(slbi_MEM), .compareS(compareS_m), .btr_cntl(btr_m), .aluOut({
        \aluOutMEM<15> , \aluOutMEM<14> , \aluOutMEM<13> , \aluOutMEM<12> , 
        \aluOutMEM<11> , \aluOutMEM<10> , \aluOutMEM<9> , \aluOutMEM<8> , 
        \aluOutMEM<7> , \aluOutMEM<6> , \aluOutMEM<5> , \aluOutMEM<4> , 
        \aluOutMEM<3> , \aluOutMEM<2> , \aluOutMEM<1> , \aluOutMEM<0> }), 
        .mem_out({\mem_out<15> , \mem_out<14> , \mem_out<13> , \mem_out<12> , 
        \mem_out<11> , \mem_out<10> , \mem_out<9> , \mem_out<8> , \mem_out<7> , 
        \mem_out<6> , \mem_out<5> , \mem_out<4> , \mem_out<3> , \mem_out<2> , 
        \mem_out<1> , \mem_out<0> }), .alu_out({\aluOutMEM<15> , 
        \aluOutMEM<14> , \aluOutMEM<13> , \aluOutMEM<12> , \aluOutMEM<11> , 
        \aluOutMEM<10> , \aluOutMEM<9> , \aluOutMEM<8> , \aluOutMEM<7> , 
        \aluOutMEM<6> , \aluOutMEM<5> , \aluOutMEM<4> , \aluOutMEM<3> , 
        \aluOutMEM<2> , \aluOutMEM<1> , \aluOutMEM<0> }), .imm({\immMEM<15> , 
        \immMEM<14> , \immMEM<13> , \immMEM<12> , \immMEM<11> , \immMEM<10> , 
        \immMEM<9> , \immMEM<8> , \immMEM<7> , \immMEM<6> , \immMEM<5> , 
        \immMEM<4> , \immMEM<3> , \immMEM<2> , \immMEM<1> , \immMEM<0> }), 
        .writereg(), .ofl(oflMEM), .zero(zeroMEM), .N(NMEM), .P(PMEM), .cout(
        c_outMEM), .inst({n952, n917, n928, n895, n941, \instMEM_normal<10> , 
        \instMEM_normal<9> , \instMEM_normal<8> , \instMEM_normal<7> , 
        \instMEM_normal<6> , \instMEM_normal<5> , \instMEM_normal<4> , 
        \instMEM_normal<3> , \instMEM_normal<2> , \instMEM_normal<1> , 
        \instMEM_normal<0> }), .ld_imm(ld_imm_m), .regwritedata({
        \regwritedata_m<15> , \regwritedata_m<14> , \regwritedata_m<13> , 
        \regwritedata_m<12> , \regwritedata_m<11> , \regwritedata_m<10> , 
        \regwritedata_m<9> , \regwritedata_m<8> , \regwritedata_m<7> , 
        \regwritedata_m<6> , \regwritedata_m<5> , \regwritedata_m<4> , 
        \regwritedata_m<3> , \regwritedata_m<2> , \regwritedata_m<1> , 
        \regwritedata_m<0> }) );
  reg3_2 rdwb ( .read({\rdWB<2> , \rdWB<1> , \rdWB<0> }), .write({\rdMEM<2> , 
        \rdMEM<1> , \rdMEM<0> }), .wr_en(n988), .rst(n986), .clk(clk) );
  reg3_1 rswb ( .read({\rsWB<2> , \rsWB<1> , \rsWB<0> }), .write({\rsMEM<2> , 
        \rsMEM<1> , \rsMEM<0> }), .wr_en(n989), .rst(n986), .clk(clk) );
  reg3_0 rwrwb ( .read({\wb_r_wr<2> , \wb_r_wr<1> , \wb_r_wr<0> }), .write({
        \mem_r_wr<2> , \mem_r_wr<1> , \mem_r_wr<0> }), .wr_en(n989), .rst(n985), .clk(clk) );
  reg16_17 instwb ( .read({\instWB_normal<15> , \instWB_normal<14> , 
        \instWB_normal<13> , \instWB_normal<12> , \instWB_normal<11> , 
        \instWB_normal<10> , \instWB_normal<9> , \instWB_normal<8> , 
        \instWB_normal<7> , \instWB_normal<6> , \instWB_normal<5> , 
        \instWB_normal<4> , \instWB_normal<3> , \instWB_normal<2> , 
        \instWB_normal<1> , \instWB_normal<0> }), .write({n952, n917, n932, 
        n957, n941, \instMEM_normal<10> , \instMEM_normal<9> , 
        \instMEM_normal<8> , \instMEM_normal<7> , \instMEM_normal<6> , 
        \instMEM_normal<5> , \instMEM_normal<4> , \instMEM_normal<3> , 
        \instMEM_normal<2> , \instMEM_normal<1> , \instMEM_normal<0> }), 
        .wr_en(n988), .rst(n985), .clk(clk) );
  reg16_16 aluOutwb ( .read({\aluOutWB<15> , \aluOutWB<14> , \aluOutWB<13> , 
        \aluOutWB<12> , \aluOutWB<11> , \aluOutWB<10> , \aluOutWB<9> , 
        \aluOutWB<8> , \aluOutWB<7> , \aluOutWB<6> , \aluOutWB<5> , 
        \aluOutWB<4> , \aluOutWB<3> , \aluOutWB<2> , \aluOutWB<1> , 
        \aluOutWB<0> }), .write({\aluOutMEM<15> , \aluOutMEM<14> , 
        \aluOutMEM<13> , \aluOutMEM<12> , \aluOutMEM<11> , \aluOutMEM<10> , 
        \aluOutMEM<9> , \aluOutMEM<8> , \aluOutMEM<7> , \aluOutMEM<6> , 
        \aluOutMEM<5> , \aluOutMEM<4> , \aluOutMEM<3> , \aluOutMEM<2> , 
        \aluOutMEM<1> , \aluOutMEM<0> }), .wr_en(n988), .rst(n986), .clk(clk)
         );
  reg16_15 memoutwb ( .read({\mem_outWB<15> , \mem_outWB<14> , \mem_outWB<13> , 
        \mem_outWB<12> , \mem_outWB<11> , \mem_outWB<10> , \mem_outWB<9> , 
        \mem_outWB<8> , \mem_outWB<7> , \mem_outWB<6> , \mem_outWB<5> , 
        \mem_outWB<4> , \mem_outWB<3> , \mem_outWB<2> , \mem_outWB<1> , 
        \mem_outWB<0> }), .write({\mem_out<15> , \mem_out<14> , \mem_out<13> , 
        \mem_out<12> , \mem_out<11> , \mem_out<10> , \mem_out<9> , 
        \mem_out<8> , \mem_out<7> , \mem_out<6> , \mem_out<5> , \mem_out<4> , 
        \mem_out<3> , \mem_out<2> , \mem_out<1> , \mem_out<0> }), .wr_en(n989), 
        .rst(n985), .clk(clk) );
  reg16_14 immwb ( .read({\immWB<15> , \immWB<14> , \immWB<13> , \immWB<12> , 
        \immWB<11> , \immWB<10> , \immWB<9> , \immWB<8> , \immWB<7> , 
        \immWB<6> , \immWB<5> , \immWB<4> , \immWB<3> , \immWB<2> , \immWB<1> , 
        \immWB<0> }), .write({\immMEM<15> , \immMEM<14> , \immMEM<13> , 
        \immMEM<12> , \immMEM<11> , \immMEM<10> , \immMEM<9> , \immMEM<8> , 
        \immMEM<7> , \immMEM<6> , \immMEM<5> , \immMEM<4> , \immMEM<3> , 
        \immMEM<2> , \immMEM<1> , \immMEM<0> }), .wr_en(n989), .rst(n986), 
        .clk(clk) );
  reg16_13 read1datawb ( .read(), .write({\read1dataMEM<15> , 
        \read1dataMEM<14> , \read1dataMEM<13> , \read1dataMEM<12> , 
        \read1dataMEM<11> , \read1dataMEM<10> , \read1dataMEM<9> , 
        \read1dataMEM<8> , \read1dataMEM<7> , \read1dataMEM<6> , 
        \read1dataMEM<5> , \read1dataMEM<4> , \read1dataMEM<3> , 
        \read1dataMEM<2> , \read1dataMEM<1> , \read1dataMEM<0> }), .wr_en(n988), .rst(n985), .clk(clk) );
  reg16_12 read2datawb ( .read(), .write({\read2dataMEM<15> , 
        \read2dataMEM<14> , \read2dataMEM<13> , \read2dataMEM<12> , 
        \read2dataMEM<11> , \read2dataMEM<10> , \read2dataMEM<9> , 
        \read2dataMEM<8> , \read2dataMEM<7> , \read2dataMEM<6> , 
        \read2dataMEM<5> , \read2dataMEM<4> , \read2dataMEM<3> , 
        \read2dataMEM<2> , \read2dataMEM<1> , \read2dataMEM<0> }), .wr_en(n989), .rst(n986), .clk(clk) );
  reg16_11 pc_inc_twowb ( .read({\pc_inc_two_WB<15> , \pc_inc_two_WB<14> , 
        \pc_inc_two_WB<13> , \pc_inc_two_WB<12> , \pc_inc_two_WB<11> , 
        \pc_inc_two_WB<10> , \pc_inc_two_WB<9> , \pc_inc_two_WB<8> , 
        \pc_inc_two_WB<7> , \pc_inc_two_WB<6> , \pc_inc_two_WB<5> , 
        \pc_inc_two_WB<4> , \pc_inc_two_WB<3> , \pc_inc_two_WB<2> , 
        \pc_inc_two_WB<1> , \pc_inc_two_WB<0> }), .write({\pc_inc_two_MEM<15> , 
        \pc_inc_two_MEM<14> , \pc_inc_two_MEM<13> , \pc_inc_two_MEM<12> , 
        \pc_inc_two_MEM<11> , \pc_inc_two_MEM<10> , \pc_inc_two_MEM<9> , 
        \pc_inc_two_MEM<8> , \pc_inc_two_MEM<7> , \pc_inc_two_MEM<6> , 
        \pc_inc_two_MEM<5> , \pc_inc_two_MEM<4> , \pc_inc_two_MEM<3> , 
        \pc_inc_two_MEM<2> , \pc_inc_two_MEM<1> , \pc_inc_two_MEM<0> }), 
        .wr_en(n988), .rst(n985), .clk(clk) );
  reg1_6 oflwb ( .d(oflMEM), .q(oflWB), .clk(clk), .rst(n986), .en(n988) );
  reg1_5 zerowb ( .d(zeroMEM), .q(zeroWB), .clk(clk), .rst(n985), .en(n1007)
         );
  reg1_4 Nwb ( .d(NMEM), .q(NWB), .clk(clk), .rst(n986), .en(n989) );
  reg1_3 Pwb ( .d(PMEM), .q(PWB), .clk(clk), .rst(n985), .en(n1007) );
  reg1_2 c_out_WB ( .d(c_outMEM), .q(c_outWB), .clk(clk), .rst(n986), .en(n989) );
  reg1_1 haltwb ( .d(haltMEM), .q(), .clk(clk), .rst(n985), .en(n1007) );
  reg1_0 slbiwb ( .d(slbi_MEM), .q(slbi_WB), .clk(clk), .rst(n986), .en(n988)
         );
  reg16_10 nx_pcwb ( .read(), .write({\nx_pcMEM<15> , \nx_pcMEM<14> , 
        \nx_pcMEM<13> , \nx_pcMEM<12> , \nx_pcMEM<11> , \nx_pcMEM<10> , 
        \nx_pcMEM<9> , \nx_pcMEM<8> , \nx_pcMEM<7> , \nx_pcMEM<6> , 
        \nx_pcMEM<5> , \nx_pcMEM<4> , \nx_pcMEM<3> , \nx_pcMEM<2> , 
        \nx_pcMEM<1> , \nx_pcMEM<0> }), .wr_en(n988), .rst(n986), .clk(clk) );
  WB_control_0 wbcntl ( .MemtoReg(memtoreg), .RegWrite(regwrite), .ld_imm(
        ld_imm), .compareS(compareS), .btr(btr), .writeR7(writeR7), .RegDst(
        regdst), .opcode({\instWB_normal<15> , \instWB_normal<14> , 
        \instWB_normal<13> , \instWB_normal<12> , \instWB_normal<11> }) );
  writeback wback ( .nxt_pc({\pc_inc_two_WB<15> , \pc_inc_two_WB<14> , 
        \pc_inc_two_WB<13> , \pc_inc_two_WB<12> , \pc_inc_two_WB<11> , 
        \pc_inc_two_WB<10> , \pc_inc_two_WB<9> , \pc_inc_two_WB<8> , 
        \pc_inc_two_WB<7> , \pc_inc_two_WB<6> , \pc_inc_two_WB<5> , 
        \pc_inc_two_WB<4> , \pc_inc_two_WB<3> , \pc_inc_two_WB<2> , 
        \pc_inc_two_WB<1> , \pc_inc_two_WB<0> }), .wr_r7(writeR7), .rd({
        \rdWB<2> , \rdWB<1> , \rdWB<0> }), .rs({\rsWB<2> , \rsWB<1> , 
        \rsWB<0> }), .regdst(regdst), .memtoreg(memtoreg), .slbi(slbi_WB), 
        .compareS(compareS), .btr_cntl(btr), .aluOut({\aluOutWB<15> , 
        \aluOutWB<14> , \aluOutWB<13> , \aluOutWB<12> , \aluOutWB<11> , 
        \aluOutWB<10> , \aluOutWB<9> , \aluOutWB<8> , \aluOutWB<7> , 
        \aluOutWB<6> , \aluOutWB<5> , \aluOutWB<4> , \aluOutWB<3> , 
        \aluOutWB<2> , \aluOutWB<1> , \aluOutWB<0> }), .mem_out({
        \mem_outWB<15> , \mem_outWB<14> , \mem_outWB<13> , \mem_outWB<12> , 
        \mem_outWB<11> , \mem_outWB<10> , \mem_outWB<9> , \mem_outWB<8> , 
        \mem_outWB<7> , \mem_outWB<6> , \mem_outWB<5> , \mem_outWB<4> , 
        \mem_outWB<3> , \mem_outWB<2> , \mem_outWB<1> , \mem_outWB<0> }), 
        .alu_out({\aluOutWB<15> , \aluOutWB<14> , \aluOutWB<13> , 
        \aluOutWB<12> , \aluOutWB<11> , \aluOutWB<10> , \aluOutWB<9> , 
        \aluOutWB<8> , \aluOutWB<7> , \aluOutWB<6> , \aluOutWB<5> , 
        \aluOutWB<4> , \aluOutWB<3> , \aluOutWB<2> , \aluOutWB<1> , 
        \aluOutWB<0> }), .imm({\immWB<15> , \immWB<14> , \immWB<13> , 
        \immWB<12> , \immWB<11> , \immWB<10> , \immWB<9> , \immWB<8> , 
        \immWB<7> , \immWB<6> , \immWB<5> , \immWB<4> , \immWB<3> , \immWB<2> , 
        \immWB<1> , \immWB<0> }), .writereg(), .ofl(oflWB), .zero(zeroWB), .N(
        NWB), .P(PWB), .cout(c_outWB), .inst({n927, n951, n949, n943, 
        \instWB_normal<11> , \instWB_normal<10> , \instWB_normal<9> , 
        \instWB_normal<8> , \instWB_normal<7> , \instWB_normal<6> , 
        \instWB_normal<5> , \instWB_normal<4> , \instWB_normal<3> , 
        \instWB_normal<2> , \instWB_normal<1> , \instWB_normal<0> }), .ld_imm(
        ld_imm), .regwritedata({\regwritedata<15> , \regwritedata<14> , 
        \regwritedata<13> , \regwritedata<12> , \regwritedata<11> , 
        \regwritedata<10> , \regwritedata<9> , \regwritedata<8> , 
        \regwritedata<7> , \regwritedata<6> , \regwritedata<5> , 
        \regwritedata<4> , \regwritedata<3> , \regwritedata<2> , 
        \regwritedata<1> , \regwritedata<0> }) );
  Harzard HDU ( .ID_rs({\r1_reg<2> , \r1_reg<1> , \r1_reg<0> }), .ID_rt({
        \r2_reg<2> , \r2_reg<1> , \r2_reg<0> }), .EX_rd({\ex_r_wr<2> , 
        \ex_r_wr<1> , \ex_r_wr<0> }), .MEM_rd({\mem_r_wr<2> , \mem_r_wr<1> , 
        \mem_r_wr<0> }), .ID_rs_v(id_rs_v), .ID_rt_v(id_rt_v), .EX_rd_v(
        ex_rd_v), .MEM_rd_v(mem_rd_v), .EX_inst({n194, n218, n181, n198, n226, 
        \instEX_normal<10> , \instEX_normal<9> , \instEX_normal<8> , 
        \instEX_normal<7> , \instEX_normal<6> , \instEX_normal<5> , 
        \instEX_normal<4> , \instEX_normal<3> , \instEX_normal<2> , 
        \instEX_normal<1> , \instEX_normal<0> }), .MEM_inst({
        \instMEM_normal<15> , n917, n932, n957, n941, \instMEM_normal<10> , 
        \instMEM_normal<9> , \instMEM_normal<8> , \instMEM_normal<7> , 
        \instMEM_normal<6> , \instMEM_normal<5> , \instMEM_normal<4> , 
        \instMEM_normal<3> , \instMEM_normal<2> , \instMEM_normal<1> , 
        \instMEM_normal<0> }), .fow_EXID_rs(fow_EXID_rs_ID), .fow_EXID_rt(
        fow_EXID_rt_ID), .fow_MEMID_rs(fow_MEMID_rs_ID), .fow_MEMID_rt(
        fow_MEMID_rt_ID), .memStall(memStall), .memDone(memDone), .memwrite(
        n796), .memread(memread), .stall(stall), .instMemStall(instMemStall), 
        .instMemDone(instMemDone), .instMemDone_q(instMemDone_q), .clk(clk), 
        .rst(n986) );
  AOI21X1 U302 ( .A(n1204), .B(n1203), .C(n989), .Y(instMemDone_d) );
  NOR3X1 U320 ( .A(jump_EX), .B(jump_ID), .C(instMemDone_q), .Y(n124) );
  INVX1 I_7 ( .A(instMemDone_q), .Y(_3_net_) );
  INVX1 U389 ( .A(n225), .Y(n177) );
  INVX4 U390 ( .A(n239), .Y(n240) );
  AND2X2 U391 ( .A(\regwritedata<13> ), .B(n1179), .Y(n547) );
  INVX2 U392 ( .A(n1007), .Y(n987) );
  INVX8 U393 ( .A(stall), .Y(n1007) );
  INVX4 U394 ( .A(n227), .Y(n872) );
  OR2X2 U395 ( .A(n1204), .B(n1003), .Y(n274) );
  INVX4 U396 ( .A(n274), .Y(n890) );
  INVX4 U397 ( .A(n632), .Y(n633) );
  INVX1 U398 ( .A(\immEX<12> ), .Y(n1039) );
  INVX1 U399 ( .A(\immEX<1> ), .Y(n1009) );
  INVX1 U400 ( .A(fow_EXID_rs_EX), .Y(n1048) );
  INVX1 U401 ( .A(n971), .Y(n899) );
  INVX1 U402 ( .A(\immEX<15> ), .Y(n1046) );
  INVX1 U403 ( .A(n864), .Y(n1196) );
  INVX1 U404 ( .A(\regwritedata_m<12> ), .Y(n1038) );
  INVX1 U405 ( .A(\rd<0> ), .Y(n1171) );
  INVX1 U406 ( .A(\rd<1> ), .Y(n1172) );
  INVX1 U407 ( .A(\rd<2> ), .Y(n1173) );
  INVX1 U408 ( .A(\rs<0> ), .Y(n1168) );
  INVX1 U409 ( .A(\rs<1> ), .Y(n1169) );
  INVX1 U410 ( .A(\rs<2> ), .Y(n1170) );
  INVX1 U411 ( .A(\instID<0> ), .Y(n1149) );
  INVX1 U412 ( .A(\instID<1> ), .Y(n1150) );
  INVX1 U413 ( .A(\instID<2> ), .Y(n1151) );
  INVX1 U414 ( .A(\instID<3> ), .Y(n1152) );
  INVX1 U415 ( .A(\instID<4> ), .Y(n1153) );
  INVX1 U416 ( .A(\instID<5> ), .Y(n1154) );
  INVX1 U417 ( .A(\instID<6> ), .Y(n1155) );
  INVX1 U418 ( .A(\instID<7> ), .Y(n1156) );
  INVX1 U419 ( .A(\instID<8> ), .Y(n1157) );
  INVX1 U420 ( .A(\instID<9> ), .Y(n1158) );
  INVX1 U421 ( .A(\instID<10> ), .Y(n1159) );
  INVX1 U422 ( .A(\instID<11> ), .Y(n1160) );
  INVX1 U423 ( .A(\instID<13> ), .Y(n1162) );
  INVX1 U424 ( .A(\instID<14> ), .Y(n1163) );
  INVX1 U425 ( .A(\instID<15> ), .Y(n1164) );
  INVX1 U426 ( .A(\immID<0> ), .Y(n1108) );
  INVX1 U427 ( .A(\immID<1> ), .Y(n1109) );
  INVX1 U428 ( .A(\immID<2> ), .Y(n1110) );
  INVX1 U429 ( .A(\immID<3> ), .Y(n1111) );
  INVX1 U430 ( .A(\immID<4> ), .Y(n1112) );
  INVX1 U431 ( .A(\immID<5> ), .Y(n1113) );
  INVX1 U432 ( .A(\immID<6> ), .Y(n1114) );
  INVX1 U433 ( .A(\displacementID<0> ), .Y(n1097) );
  INVX1 U434 ( .A(\displacementID<1> ), .Y(n1098) );
  INVX1 U435 ( .A(\displacementID<2> ), .Y(n1099) );
  INVX1 U436 ( .A(\displacementID<3> ), .Y(n1100) );
  INVX1 U437 ( .A(\displacementID<4> ), .Y(n1101) );
  INVX1 U438 ( .A(\displacementID<5> ), .Y(n1102) );
  INVX1 U439 ( .A(\displacementID<6> ), .Y(n1103) );
  INVX1 U440 ( .A(\displacementID<7> ), .Y(n1104) );
  INVX1 U441 ( .A(\displacementID<8> ), .Y(n1105) );
  INVX1 U442 ( .A(\displacementID<9> ), .Y(n1106) );
  INVX1 U443 ( .A(\displacementID<10> ), .Y(n1107) );
  INVX1 U444 ( .A(haltID), .Y(n1095) );
  INVX1 U445 ( .A(\pc_inc_two_ID<0> ), .Y(n1079) );
  INVX1 U446 ( .A(\pc_inc_two_ID<1> ), .Y(n1080) );
  INVX1 U447 ( .A(\pc_inc_two_ID<2> ), .Y(n1081) );
  INVX1 U448 ( .A(\pc_inc_two_ID<3> ), .Y(n1082) );
  INVX1 U449 ( .A(\pc_inc_two_ID<4> ), .Y(n1083) );
  INVX1 U450 ( .A(\pc_inc_two_ID<5> ), .Y(n1084) );
  INVX1 U451 ( .A(\pc_inc_two_ID<6> ), .Y(n1085) );
  INVX1 U452 ( .A(\pc_inc_two_ID<7> ), .Y(n1086) );
  INVX1 U453 ( .A(\pc_inc_two_ID<8> ), .Y(n1087) );
  INVX1 U454 ( .A(\pc_inc_two_ID<9> ), .Y(n1088) );
  INVX1 U455 ( .A(\pc_inc_two_ID<10> ), .Y(n1089) );
  INVX1 U456 ( .A(\pc_inc_two_ID<11> ), .Y(n1090) );
  INVX1 U457 ( .A(\pc_inc_two_ID<12> ), .Y(n1091) );
  INVX1 U458 ( .A(\pc_inc_two_ID<13> ), .Y(n1092) );
  INVX1 U459 ( .A(\pc_inc_two_ID<14> ), .Y(n1093) );
  INVX1 U460 ( .A(\pc_inc_two_ID<15> ), .Y(n1094) );
  INVX1 U461 ( .A(fow_EXID_rs_ID), .Y(n1078) );
  INVX1 U462 ( .A(fow_MEMID_rs_ID), .Y(n1077) );
  INVX1 U463 ( .A(fow_EXID_rt_ID), .Y(n1076) );
  INVX1 U464 ( .A(fow_MEMID_rt_ID), .Y(n1075) );
  INVX1 U465 ( .A(jmp_r_ID), .Y(n1074) );
  INVX1 U466 ( .A(\nx_pcID<0> ), .Y(n1058) );
  INVX1 U467 ( .A(\nx_pcID<1> ), .Y(n1059) );
  INVX1 U468 ( .A(\nx_pcID<2> ), .Y(n1060) );
  INVX1 U469 ( .A(\nx_pcID<3> ), .Y(n1061) );
  INVX1 U470 ( .A(\nx_pcID<4> ), .Y(n1062) );
  INVX1 U471 ( .A(\nx_pcID<5> ), .Y(n1063) );
  INVX1 U472 ( .A(\nx_pcID<6> ), .Y(n1064) );
  INVX1 U473 ( .A(\nx_pcID<7> ), .Y(n1065) );
  INVX1 U474 ( .A(\nx_pcID<8> ), .Y(n1066) );
  INVX1 U475 ( .A(\nx_pcID<9> ), .Y(n1067) );
  INVX1 U476 ( .A(\nx_pcID<10> ), .Y(n1068) );
  INVX1 U477 ( .A(\nx_pcID<11> ), .Y(n1069) );
  INVX1 U478 ( .A(\nx_pcID<12> ), .Y(n1070) );
  INVX1 U479 ( .A(\nx_pcID<13> ), .Y(n1071) );
  INVX1 U480 ( .A(\nx_pcID<14> ), .Y(n1072) );
  INVX1 U481 ( .A(\nx_pcID<15> ), .Y(n1073) );
  INVX1 U482 ( .A(branch_id), .Y(n1057) );
  AND2X1 U483 ( .A(n859), .B(n703), .Y(n760) );
  AND2X1 U484 ( .A(n229), .B(n564), .Y(n219) );
  INVX1 U485 ( .A(n863), .Y(n1020) );
  BUFX2 U486 ( .A(n124), .Y(n991) );
  INVX1 U487 ( .A(instMemDone), .Y(n1203) );
  AND2X1 U488 ( .A(n1200), .B(n858), .Y(n753) );
  INVX1 U489 ( .A(n1197), .Y(n209) );
  INVX1 U490 ( .A(n835), .Y(n1188) );
  INVX2 U491 ( .A(n638), .Y(n639) );
  INVX2 U492 ( .A(n967), .Y(\opB<10> ) );
  INVX1 U493 ( .A(n235), .Y(n236) );
  INVX1 U494 ( .A(jump_EX), .Y(n1175) );
  INVX1 U495 ( .A(\instID<12> ), .Y(n1161) );
  AND2X1 U496 ( .A(n179), .B(n701), .Y(n782) );
  AND2X1 U497 ( .A(n694), .B(n700), .Y(n780) );
  AND2X1 U498 ( .A(n692), .B(n858), .Y(n778) );
  AND2X1 U499 ( .A(n690), .B(n699), .Y(n772) );
  AND2X1 U500 ( .A(n688), .B(n698), .Y(n770) );
  AND2X1 U501 ( .A(n686), .B(n697), .Y(n768) );
  AND2X1 U502 ( .A(n1187), .B(n707), .Y(n766) );
  AND2X1 U503 ( .A(n1186), .B(n705), .Y(n764) );
  INVX8 U504 ( .A(n883), .Y(n998) );
  INVX8 U505 ( .A(n1053), .Y(n1056) );
  AND2X2 U506 ( .A(fow_EXID_rt_EX), .B(n191), .Y(n178) );
  INVX4 U507 ( .A(n994), .Y(n1006) );
  INVX8 U508 ( .A(n884), .Y(n1002) );
  INVX1 U509 ( .A(\immID<13> ), .Y(n1116) );
  INVX1 U510 ( .A(n841), .Y(n179) );
  INVX4 U511 ( .A(n634), .Y(n243) );
  BUFX2 U512 ( .A(\regwritedata_m<10> ), .Y(n180) );
  BUFX2 U513 ( .A(\instEX_normal<13> ), .Y(n181) );
  INVX1 U514 ( .A(n921), .Y(n182) );
  INVX2 U515 ( .A(n220), .Y(n873) );
  AND2X2 U516 ( .A(\regwritedata<10> ), .B(n285), .Y(n969) );
  INVX1 U517 ( .A(n276), .Y(n211) );
  AND2X1 U518 ( .A(\regwritedata_m<7> ), .B(n178), .Y(n662) );
  INVX1 U519 ( .A(\regwritedata_m<5> ), .Y(n183) );
  INVX1 U520 ( .A(n183), .Y(n184) );
  BUFX2 U521 ( .A(n295), .Y(n185) );
  AND2X2 U522 ( .A(n922), .B(n923), .Y(n186) );
  INVX2 U523 ( .A(n294), .Y(n295) );
  BUFX2 U524 ( .A(n718), .Y(n187) );
  AND2X2 U525 ( .A(\regwritedata_m<4> ), .B(fow_EXID_rs_EX), .Y(n1050) );
  INVX8 U526 ( .A(n984), .Y(\forwarded_read1dataEX<5> ) );
  OR2X2 U527 ( .A(n306), .B(n719), .Y(n188) );
  INVX1 U528 ( .A(n880), .Y(n189) );
  INVX1 U529 ( .A(alusrc), .Y(n190) );
  INVX4 U530 ( .A(n190), .Y(n191) );
  INVX1 U531 ( .A(alusrc), .Y(n192) );
  INVX1 U532 ( .A(n192), .Y(n193) );
  AND2X2 U533 ( .A(n191), .B(n744), .Y(n722) );
  BUFX2 U534 ( .A(\instEX_normal<15> ), .Y(n194) );
  INVX1 U535 ( .A(\regwritedata_m<0> ), .Y(n195) );
  INVX1 U536 ( .A(n195), .Y(n196) );
  INVX1 U537 ( .A(n203), .Y(n197) );
  BUFX2 U538 ( .A(n236), .Y(n198) );
  INVX1 U539 ( .A(n191), .Y(n208) );
  INVX4 U540 ( .A(n193), .Y(n1036) );
  INVX1 U541 ( .A(\regwritedata_m<0> ), .Y(n199) );
  BUFX2 U542 ( .A(\forwarded_read1dataEX<8> ), .Y(n200) );
  NOR3X1 U543 ( .A(n202), .B(n296), .C(n787), .Y(n201) );
  INVX2 U544 ( .A(n201), .Y(\opB<13> ) );
  INVX1 U545 ( .A(n1040), .Y(n202) );
  INVX1 U546 ( .A(\regwritedata<7> ), .Y(n203) );
  AND2X2 U547 ( .A(\regwritedata_m<13> ), .B(fow_EXID_rt_EX), .Y(n569) );
  BUFX2 U548 ( .A(n177), .Y(n204) );
  BUFX2 U549 ( .A(\opB<2> ), .Y(n205) );
  AND2X1 U550 ( .A(\regwritedata_m<14> ), .B(fow_EXID_rt_EX), .Y(n603) );
  OR2X2 U551 ( .A(n981), .B(n659), .Y(n206) );
  INVX2 U552 ( .A(n904), .Y(\forwarded_read1dataEX<8> ) );
  AND2X2 U553 ( .A(\regwritedata<3> ), .B(n285), .Y(n290) );
  NOR3X1 U554 ( .A(n208), .B(n209), .C(n210), .Y(n207) );
  INVX1 U555 ( .A(\regwritedata<8> ), .Y(n210) );
  AND2X2 U556 ( .A(n292), .B(n643), .Y(n762) );
  INVX4 U557 ( .A(n961), .Y(n962) );
  AND2X2 U558 ( .A(\regwritedata_m<10> ), .B(n1032), .Y(n679) );
  AND2X2 U559 ( .A(n180), .B(fow_EXID_rt_EX), .Y(n687) );
  BUFX2 U560 ( .A(\regwritedata<8> ), .Y(n212) );
  OR2X2 U561 ( .A(n290), .B(n214), .Y(n213) );
  INVX1 U562 ( .A(n1023), .Y(n214) );
  INVX1 U563 ( .A(n654), .Y(n215) );
  AND2X2 U564 ( .A(n310), .B(n840), .Y(n673) );
  INVX1 U565 ( .A(n283), .Y(n216) );
  BUFX2 U566 ( .A(\regwritedata<13> ), .Y(n217) );
  AND2X2 U567 ( .A(\immEX<4> ), .B(n925), .Y(n710) );
  INVX1 U568 ( .A(n925), .Y(n1047) );
  AND2X2 U569 ( .A(\immEX<9> ), .B(n925), .Y(n714) );
  BUFX2 U570 ( .A(\instEX_normal<14> ), .Y(n218) );
  NOR3X1 U571 ( .A(n738), .B(n298), .C(n788), .Y(n220) );
  INVX1 U572 ( .A(n913), .Y(n221) );
  INVX1 U573 ( .A(n221), .Y(n222) );
  OR2X2 U574 ( .A(n547), .B(n674), .Y(n223) );
  AND2X2 U575 ( .A(n217), .B(n1197), .Y(n706) );
  INVX1 U576 ( .A(n901), .Y(n224) );
  INVX1 U577 ( .A(\regwritedata<1> ), .Y(n225) );
  INVX1 U578 ( .A(n204), .Y(n1200) );
  AND2X2 U579 ( .A(n204), .B(n1197), .Y(n691) );
  AND2X2 U580 ( .A(\immEX<6> ), .B(n186), .Y(n712) );
  AND2X2 U581 ( .A(n923), .B(n924), .Y(n784) );
  BUFX2 U582 ( .A(\instEX_normal<11> ), .Y(n226) );
  AND2X2 U583 ( .A(\regwritedata<2> ), .B(n1179), .Y(n605) );
  INVX1 U584 ( .A(n191), .Y(n1019) );
  NOR3X1 U585 ( .A(n786), .B(n293), .C(n207), .Y(n227) );
  AND2X2 U586 ( .A(n275), .B(n187), .Y(n671) );
  OR2X2 U587 ( .A(n550), .B(n232), .Y(n228) );
  INVX1 U588 ( .A(n233), .Y(n1027) );
  INVX1 U589 ( .A(n1011), .Y(n230) );
  NOR3X1 U590 ( .A(n878), .B(n865), .C(n230), .Y(n229) );
  INVX1 U591 ( .A(n970), .Y(\forwarded_read1dataEX<15> ) );
  INVX1 U592 ( .A(n970), .Y(n882) );
  BUFX2 U593 ( .A(\regwritedata<2> ), .Y(n231) );
  AND2X2 U594 ( .A(n1013), .B(n566), .Y(n615) );
  OAI21X1 U595 ( .A(n678), .B(n199), .C(n281), .Y(n232) );
  BUFX2 U596 ( .A(\regwritedata<11> ), .Y(n909) );
  NOR3X1 U597 ( .A(n833), .B(n850), .C(n651), .Y(n233) );
  INVX1 U598 ( .A(n543), .Y(n868) );
  AND2X2 U599 ( .A(\regwritedata_m<4> ), .B(fow_EXID_rt_EX), .Y(n851) );
  INVX4 U600 ( .A(n936), .Y(\opB<2> ) );
  NOR3X1 U601 ( .A(n867), .B(n307), .C(n621), .Y(n234) );
  INVX2 U602 ( .A(n234), .Y(n902) );
  INVX2 U603 ( .A(n282), .Y(n870) );
  INVX1 U604 ( .A(\instEX_normal<12> ), .Y(n235) );
  AND2X2 U605 ( .A(n275), .B(n718), .Y(n237) );
  INVX1 U606 ( .A(n237), .Y(n238) );
  AND2X2 U607 ( .A(n215), .B(n592), .Y(n239) );
  AND2X2 U608 ( .A(n642), .B(n292), .Y(n241) );
  INVX1 U609 ( .A(n241), .Y(n242) );
  OR2X2 U610 ( .A(n1002), .B(n1183), .Y(n244) );
  INVX1 U611 ( .A(n244), .Y(n245) );
  OR2X2 U612 ( .A(n1002), .B(n1057), .Y(n246) );
  INVX1 U613 ( .A(n246), .Y(n247) );
  OR2X2 U614 ( .A(n1002), .B(n1058), .Y(n248) );
  INVX1 U615 ( .A(n248), .Y(n249) );
  OR2X2 U616 ( .A(n1002), .B(n1060), .Y(n250) );
  INVX1 U617 ( .A(n250), .Y(n251) );
  OR2X2 U618 ( .A(n1002), .B(n1062), .Y(n252) );
  INVX1 U619 ( .A(n252), .Y(n253) );
  OR2X2 U620 ( .A(n1002), .B(n1064), .Y(n254) );
  INVX1 U621 ( .A(n254), .Y(n255) );
  OR2X2 U622 ( .A(n1002), .B(n1066), .Y(n256) );
  INVX1 U623 ( .A(n256), .Y(n257) );
  OR2X2 U624 ( .A(n1002), .B(n1068), .Y(n258) );
  INVX1 U625 ( .A(n258), .Y(n259) );
  OR2X2 U626 ( .A(n1002), .B(n1070), .Y(n260) );
  INVX1 U627 ( .A(n260), .Y(n261) );
  OR2X2 U628 ( .A(n1002), .B(n1072), .Y(n262) );
  INVX1 U629 ( .A(n262), .Y(n263) );
  OR2X2 U630 ( .A(n1002), .B(n1075), .Y(n264) );
  INVX1 U631 ( .A(n264), .Y(n265) );
  OR2X2 U632 ( .A(n1002), .B(n1078), .Y(n266) );
  INVX1 U633 ( .A(n266), .Y(n267) );
  OR2X2 U634 ( .A(n1002), .B(n1079), .Y(n268) );
  INVX1 U635 ( .A(n268), .Y(n269) );
  OR2X2 U636 ( .A(n1002), .B(n1081), .Y(n270) );
  INVX1 U637 ( .A(n270), .Y(n271) );
  OR2X2 U638 ( .A(n997), .B(n1161), .Y(n272) );
  INVX1 U639 ( .A(n272), .Y(n273) );
  AND2X2 U640 ( .A(n723), .B(n663), .Y(n275) );
  AND2X2 U641 ( .A(n596), .B(n279), .Y(n276) );
  INVX1 U642 ( .A(n276), .Y(n277) );
  AND2X2 U643 ( .A(\regwritedata<11> ), .B(n1179), .Y(n278) );
  INVX1 U644 ( .A(n278), .Y(n279) );
  AND2X2 U645 ( .A(n287), .B(n598), .Y(n280) );
  AND2X2 U646 ( .A(n280), .B(n600), .Y(n281) );
  AND2X2 U647 ( .A(n609), .B(n590), .Y(n282) );
  AND2X2 U648 ( .A(n721), .B(n589), .Y(n283) );
  INVX1 U649 ( .A(n283), .Y(n284) );
  AND2X2 U650 ( .A(n191), .B(n1197), .Y(n285) );
  AND2X2 U651 ( .A(n191), .B(n743), .Y(n286) );
  INVX1 U652 ( .A(n286), .Y(n287) );
  AND2X2 U653 ( .A(n191), .B(n602), .Y(n288) );
  INVX1 U654 ( .A(n288), .Y(n289) );
  AND2X2 U655 ( .A(n285), .B(n667), .Y(n291) );
  INVX1 U656 ( .A(n291), .Y(n292) );
  AND2X2 U657 ( .A(n645), .B(n191), .Y(n293) );
  AND2X2 U658 ( .A(n591), .B(n611), .Y(n294) );
  AND2X2 U659 ( .A(n191), .B(n648), .Y(n296) );
  AND2X2 U660 ( .A(n729), .B(n604), .Y(n297) );
  AND2X2 U661 ( .A(n191), .B(n797), .Y(n298) );
  AND2X2 U662 ( .A(n191), .B(\forwarded_read2dataEX<15> ), .Y(n299) );
  INVX1 U663 ( .A(n299), .Y(n300) );
  AND2X2 U664 ( .A(n655), .B(n594), .Y(n301) );
  AND2X2 U665 ( .A(n613), .B(n650), .Y(n302) );
  INVX1 U666 ( .A(n302), .Y(n303) );
  AND2X2 U667 ( .A(\regwritedata<3> ), .B(n1179), .Y(n304) );
  INVX1 U668 ( .A(n304), .Y(n305) );
  AND2X2 U669 ( .A(n1179), .B(n911), .Y(n306) );
  AND2X2 U670 ( .A(\regwritedata_m<9> ), .B(fow_EXID_rs_EX), .Y(n307) );
  AND2X2 U671 ( .A(fow_EXID_rs_EX), .B(\regwritedata_m<11> ), .Y(n308) );
  AND2X2 U672 ( .A(fow_EXID_rs_EX), .B(\regwritedata_m<13> ), .Y(n309) );
  INVX1 U673 ( .A(n309), .Y(n310) );
  OR2X2 U674 ( .A(n998), .B(n1059), .Y(n311) );
  INVX1 U675 ( .A(n311), .Y(n312) );
  OR2X2 U676 ( .A(n998), .B(n1061), .Y(n313) );
  INVX1 U677 ( .A(n313), .Y(n314) );
  OR2X2 U678 ( .A(n998), .B(n1063), .Y(n315) );
  INVX1 U679 ( .A(n315), .Y(n316) );
  OR2X2 U680 ( .A(n998), .B(n1065), .Y(n317) );
  INVX1 U681 ( .A(n317), .Y(n318) );
  OR2X2 U682 ( .A(n998), .B(n1067), .Y(n319) );
  INVX1 U683 ( .A(n319), .Y(n320) );
  OR2X2 U684 ( .A(n998), .B(n1069), .Y(n321) );
  INVX1 U685 ( .A(n321), .Y(n322) );
  OR2X2 U686 ( .A(n997), .B(n1071), .Y(n323) );
  INVX1 U687 ( .A(n323), .Y(n324) );
  OR2X2 U688 ( .A(n996), .B(n1073), .Y(n325) );
  INVX1 U689 ( .A(n325), .Y(n326) );
  OR2X1 U690 ( .A(n996), .B(n1074), .Y(n327) );
  INVX1 U691 ( .A(n327), .Y(n328) );
  OR2X1 U692 ( .A(n998), .B(n1076), .Y(n329) );
  INVX1 U693 ( .A(n329), .Y(n330) );
  OR2X1 U694 ( .A(n997), .B(n1077), .Y(n331) );
  INVX1 U695 ( .A(n331), .Y(n332) );
  OR2X1 U696 ( .A(n998), .B(n1080), .Y(n333) );
  INVX1 U697 ( .A(n333), .Y(n334) );
  OR2X1 U698 ( .A(n996), .B(n1082), .Y(n335) );
  INVX1 U699 ( .A(n335), .Y(n336) );
  OR2X2 U700 ( .A(n999), .B(n1083), .Y(n337) );
  INVX1 U701 ( .A(n337), .Y(n338) );
  OR2X2 U702 ( .A(n885), .B(n1084), .Y(n339) );
  INVX1 U703 ( .A(n339), .Y(n340) );
  OR2X2 U704 ( .A(n885), .B(n1085), .Y(n341) );
  INVX1 U705 ( .A(n341), .Y(n342) );
  OR2X2 U706 ( .A(n999), .B(n1086), .Y(n343) );
  INVX1 U707 ( .A(n343), .Y(n344) );
  OR2X2 U708 ( .A(n1001), .B(n1087), .Y(n345) );
  INVX1 U709 ( .A(n345), .Y(n346) );
  OR2X2 U710 ( .A(n1000), .B(n1088), .Y(n347) );
  INVX1 U711 ( .A(n347), .Y(n348) );
  OR2X2 U712 ( .A(n885), .B(n1089), .Y(n349) );
  INVX1 U713 ( .A(n349), .Y(n350) );
  OR2X2 U714 ( .A(n885), .B(n1090), .Y(n351) );
  INVX1 U715 ( .A(n351), .Y(n352) );
  OR2X2 U716 ( .A(n1001), .B(n1091), .Y(n353) );
  INVX1 U717 ( .A(n353), .Y(n354) );
  OR2X2 U718 ( .A(n1000), .B(n1092), .Y(n355) );
  INVX1 U719 ( .A(n355), .Y(n356) );
  OR2X2 U720 ( .A(n999), .B(n1093), .Y(n357) );
  INVX1 U721 ( .A(n357), .Y(n358) );
  OR2X2 U722 ( .A(n885), .B(n1094), .Y(n359) );
  INVX1 U723 ( .A(n359), .Y(n360) );
  OR2X2 U724 ( .A(n1000), .B(n1095), .Y(n361) );
  INVX1 U725 ( .A(n361), .Y(n362) );
  OR2X2 U726 ( .A(n1000), .B(n1096), .Y(n363) );
  INVX1 U727 ( .A(n363), .Y(n364) );
  OR2X2 U728 ( .A(n999), .B(n1097), .Y(n365) );
  INVX1 U729 ( .A(n365), .Y(n366) );
  OR2X2 U730 ( .A(n1001), .B(n1098), .Y(n367) );
  INVX1 U731 ( .A(n367), .Y(n368) );
  OR2X2 U732 ( .A(n1000), .B(n1099), .Y(n369) );
  INVX1 U733 ( .A(n369), .Y(n370) );
  OR2X2 U734 ( .A(n885), .B(n1100), .Y(n371) );
  INVX1 U735 ( .A(n371), .Y(n372) );
  OR2X2 U736 ( .A(n885), .B(n1101), .Y(n373) );
  INVX1 U737 ( .A(n373), .Y(n374) );
  OR2X2 U738 ( .A(n1001), .B(n1102), .Y(n375) );
  INVX1 U739 ( .A(n375), .Y(n376) );
  OR2X2 U740 ( .A(n1000), .B(n1103), .Y(n377) );
  INVX1 U741 ( .A(n377), .Y(n378) );
  OR2X2 U742 ( .A(n999), .B(n1104), .Y(n379) );
  INVX1 U743 ( .A(n379), .Y(n380) );
  OR2X2 U744 ( .A(n885), .B(n1105), .Y(n381) );
  INVX1 U745 ( .A(n381), .Y(n382) );
  OR2X2 U746 ( .A(n885), .B(n1106), .Y(n383) );
  INVX1 U747 ( .A(n383), .Y(n384) );
  OR2X2 U748 ( .A(n1001), .B(n1107), .Y(n385) );
  INVX1 U749 ( .A(n385), .Y(n386) );
  OR2X2 U750 ( .A(n997), .B(n1108), .Y(n387) );
  INVX1 U751 ( .A(n387), .Y(n388) );
  OR2X2 U752 ( .A(n997), .B(n1109), .Y(n389) );
  INVX1 U753 ( .A(n389), .Y(n390) );
  OR2X2 U754 ( .A(n997), .B(n1110), .Y(n391) );
  INVX1 U755 ( .A(n391), .Y(n392) );
  OR2X2 U756 ( .A(n997), .B(n1111), .Y(n393) );
  INVX1 U757 ( .A(n393), .Y(n394) );
  OR2X2 U758 ( .A(n996), .B(n1112), .Y(n395) );
  INVX1 U759 ( .A(n395), .Y(n396) );
  OR2X2 U760 ( .A(n997), .B(n1113), .Y(n397) );
  INVX1 U761 ( .A(n397), .Y(n398) );
  OR2X2 U762 ( .A(n996), .B(n1114), .Y(n399) );
  INVX1 U763 ( .A(n399), .Y(n400) );
  OR2X2 U764 ( .A(n997), .B(n1115), .Y(n401) );
  INVX1 U765 ( .A(n401), .Y(n402) );
  INVX1 U766 ( .A(n404), .Y(n403) );
  OR2X2 U767 ( .A(n999), .B(n1116), .Y(n404) );
  OR2X2 U768 ( .A(n885), .B(n1117), .Y(n405) );
  INVX1 U769 ( .A(n405), .Y(n406) );
  OR2X2 U770 ( .A(n885), .B(n1118), .Y(n407) );
  INVX1 U771 ( .A(n407), .Y(n408) );
  OR2X2 U772 ( .A(n1001), .B(n1119), .Y(n409) );
  INVX1 U773 ( .A(n409), .Y(n410) );
  OR2X2 U774 ( .A(n1000), .B(n1120), .Y(n411) );
  INVX1 U775 ( .A(n411), .Y(n412) );
  OR2X2 U776 ( .A(n999), .B(n1121), .Y(n413) );
  INVX1 U777 ( .A(n413), .Y(n414) );
  OR2X2 U778 ( .A(n885), .B(n1122), .Y(n415) );
  INVX1 U779 ( .A(n415), .Y(n416) );
  OR2X2 U780 ( .A(n885), .B(n1123), .Y(n417) );
  INVX1 U781 ( .A(n417), .Y(n418) );
  OR2X2 U782 ( .A(n1001), .B(n1124), .Y(n419) );
  INVX1 U783 ( .A(n419), .Y(n420) );
  OR2X2 U784 ( .A(n1000), .B(n1125), .Y(n421) );
  INVX1 U785 ( .A(n421), .Y(n422) );
  OR2X2 U786 ( .A(n999), .B(n1126), .Y(n423) );
  INVX1 U787 ( .A(n423), .Y(n424) );
  OR2X2 U788 ( .A(n885), .B(n1127), .Y(n425) );
  INVX1 U789 ( .A(n425), .Y(n426) );
  OR2X2 U790 ( .A(n885), .B(n1128), .Y(n427) );
  INVX1 U791 ( .A(n427), .Y(n428) );
  OR2X2 U792 ( .A(n999), .B(n1129), .Y(n429) );
  INVX1 U793 ( .A(n429), .Y(n430) );
  OR2X2 U794 ( .A(n885), .B(n1130), .Y(n431) );
  INVX1 U795 ( .A(n431), .Y(n432) );
  OR2X2 U796 ( .A(n885), .B(n1131), .Y(n433) );
  INVX1 U797 ( .A(n433), .Y(n434) );
  OR2X2 U798 ( .A(n1001), .B(n1132), .Y(n435) );
  INVX1 U799 ( .A(n435), .Y(n436) );
  OR2X2 U800 ( .A(n885), .B(n1133), .Y(n437) );
  INVX1 U801 ( .A(n437), .Y(n438) );
  OR2X2 U802 ( .A(n885), .B(n1134), .Y(n439) );
  INVX1 U803 ( .A(n439), .Y(n440) );
  OR2X2 U804 ( .A(n1001), .B(n1135), .Y(n441) );
  INVX1 U805 ( .A(n441), .Y(n442) );
  OR2X1 U806 ( .A(n998), .B(n1136), .Y(n443) );
  INVX1 U807 ( .A(n443), .Y(n444) );
  OR2X1 U808 ( .A(n998), .B(n1137), .Y(n445) );
  INVX1 U809 ( .A(n445), .Y(n446) );
  OR2X1 U810 ( .A(n998), .B(n1138), .Y(n447) );
  INVX1 U811 ( .A(n447), .Y(n448) );
  OR2X1 U812 ( .A(n998), .B(n1139), .Y(n449) );
  INVX1 U813 ( .A(n449), .Y(n450) );
  OR2X1 U814 ( .A(n998), .B(n1140), .Y(n451) );
  INVX1 U815 ( .A(n451), .Y(n452) );
  OR2X1 U816 ( .A(n998), .B(n1141), .Y(n453) );
  INVX1 U817 ( .A(n453), .Y(n454) );
  OR2X1 U818 ( .A(n998), .B(n1142), .Y(n455) );
  INVX1 U819 ( .A(n455), .Y(n456) );
  OR2X1 U820 ( .A(n998), .B(n1143), .Y(n457) );
  INVX1 U821 ( .A(n457), .Y(n458) );
  OR2X1 U822 ( .A(n998), .B(n1144), .Y(n459) );
  INVX1 U823 ( .A(n459), .Y(n460) );
  OR2X1 U824 ( .A(n998), .B(n1145), .Y(n461) );
  INVX1 U825 ( .A(n461), .Y(n462) );
  OR2X1 U826 ( .A(n998), .B(n1146), .Y(n463) );
  INVX1 U827 ( .A(n463), .Y(n464) );
  OR2X1 U828 ( .A(n998), .B(n1147), .Y(n465) );
  INVX1 U829 ( .A(n465), .Y(n466) );
  OR2X1 U830 ( .A(n998), .B(n1148), .Y(n467) );
  INVX1 U831 ( .A(n467), .Y(n468) );
  OR2X2 U832 ( .A(n997), .B(n1149), .Y(n469) );
  INVX1 U833 ( .A(n469), .Y(n470) );
  OR2X2 U834 ( .A(n997), .B(n1150), .Y(n471) );
  INVX1 U835 ( .A(n471), .Y(n472) );
  OR2X2 U836 ( .A(n997), .B(n1151), .Y(n473) );
  INVX1 U837 ( .A(n473), .Y(n474) );
  OR2X2 U838 ( .A(n997), .B(n1152), .Y(n475) );
  INVX1 U839 ( .A(n475), .Y(n476) );
  OR2X2 U840 ( .A(n997), .B(n1153), .Y(n477) );
  INVX1 U841 ( .A(n477), .Y(n478) );
  OR2X2 U842 ( .A(n997), .B(n1154), .Y(n479) );
  INVX1 U843 ( .A(n479), .Y(n480) );
  OR2X2 U844 ( .A(n997), .B(n1155), .Y(n481) );
  INVX1 U845 ( .A(n481), .Y(n482) );
  OR2X2 U846 ( .A(n997), .B(n1156), .Y(n483) );
  INVX1 U847 ( .A(n483), .Y(n484) );
  OR2X2 U848 ( .A(n997), .B(n1157), .Y(n485) );
  INVX1 U849 ( .A(n485), .Y(n486) );
  OR2X2 U850 ( .A(n997), .B(n1158), .Y(n487) );
  INVX1 U851 ( .A(n487), .Y(n488) );
  OR2X2 U852 ( .A(n997), .B(n1159), .Y(n489) );
  INVX1 U853 ( .A(n489), .Y(n490) );
  OR2X2 U854 ( .A(n997), .B(n1162), .Y(n491) );
  INVX1 U855 ( .A(n491), .Y(n492) );
  OR2X2 U856 ( .A(n996), .B(n1163), .Y(n493) );
  INVX1 U857 ( .A(n493), .Y(n494) );
  OR2X2 U858 ( .A(n996), .B(n1164), .Y(n495) );
  INVX1 U859 ( .A(n495), .Y(n496) );
  OR2X2 U860 ( .A(n996), .B(n1165), .Y(n497) );
  INVX1 U861 ( .A(n497), .Y(n498) );
  OR2X2 U862 ( .A(n996), .B(n1166), .Y(n499) );
  INVX1 U863 ( .A(n499), .Y(n500) );
  OR2X2 U864 ( .A(n996), .B(n1167), .Y(n501) );
  INVX1 U865 ( .A(n501), .Y(n502) );
  OR2X2 U866 ( .A(n996), .B(n1168), .Y(n503) );
  INVX1 U867 ( .A(n503), .Y(n504) );
  OR2X2 U868 ( .A(n996), .B(n1169), .Y(n505) );
  INVX1 U869 ( .A(n505), .Y(n506) );
  OR2X2 U870 ( .A(n996), .B(n1170), .Y(n507) );
  INVX1 U871 ( .A(n507), .Y(n508) );
  OR2X2 U872 ( .A(n996), .B(n1171), .Y(n509) );
  INVX1 U873 ( .A(n509), .Y(n510) );
  OR2X2 U874 ( .A(n996), .B(n1172), .Y(n511) );
  INVX1 U875 ( .A(n511), .Y(n512) );
  OR2X2 U876 ( .A(n996), .B(n1173), .Y(n513) );
  INVX1 U877 ( .A(n513), .Y(n514) );
  OR2X2 U878 ( .A(n731), .B(n996), .Y(n515) );
  INVX1 U879 ( .A(n515), .Y(n516) );
  OR2X2 U880 ( .A(n733), .B(n996), .Y(n517) );
  INVX1 U881 ( .A(n517), .Y(n518) );
  AND2X2 U882 ( .A(\instIF_q<0> ), .B(n918), .Y(n519) );
  INVX1 U883 ( .A(n519), .Y(n520) );
  AND2X2 U884 ( .A(\instIF_q<1> ), .B(n918), .Y(n521) );
  INVX1 U885 ( .A(n521), .Y(n522) );
  AND2X2 U886 ( .A(\instIF_q<2> ), .B(n918), .Y(n523) );
  INVX1 U887 ( .A(n523), .Y(n524) );
  AND2X2 U888 ( .A(\instIF_q<3> ), .B(n918), .Y(n525) );
  INVX1 U889 ( .A(n525), .Y(n526) );
  AND2X2 U890 ( .A(\instIF_q<4> ), .B(n918), .Y(n527) );
  INVX1 U891 ( .A(n527), .Y(n528) );
  AND2X2 U892 ( .A(\instIF_q<6> ), .B(n918), .Y(n529) );
  INVX1 U893 ( .A(n529), .Y(n530) );
  AND2X2 U894 ( .A(\instIF_q<7> ), .B(n890), .Y(n531) );
  INVX1 U895 ( .A(n531), .Y(n532) );
  AND2X2 U896 ( .A(\instIF_q<8> ), .B(n918), .Y(n533) );
  INVX1 U897 ( .A(n533), .Y(n534) );
  AND2X2 U898 ( .A(\instIF_q<9> ), .B(n890), .Y(n535) );
  INVX1 U899 ( .A(n535), .Y(n536) );
  AND2X2 U900 ( .A(\instIF_q<10> ), .B(n918), .Y(n537) );
  INVX1 U901 ( .A(n537), .Y(n538) );
  AND2X2 U902 ( .A(\instIF_q<12> ), .B(n890), .Y(n539) );
  INVX1 U903 ( .A(n539), .Y(n540) );
  AND2X2 U904 ( .A(\instIF_q<13> ), .B(n918), .Y(n541) );
  INVX1 U905 ( .A(n541), .Y(n542) );
  AND2X2 U906 ( .A(n653), .B(n606), .Y(n543) );
  INVX1 U907 ( .A(n543), .Y(n544) );
  BUFX2 U908 ( .A(n1051), .Y(n545) );
  BUFX2 U909 ( .A(n1052), .Y(n546) );
  AND2X2 U910 ( .A(n1179), .B(\regwritedata<15> ), .Y(n548) );
  INVX1 U911 ( .A(n548), .Y(n549) );
  AND2X2 U912 ( .A(n285), .B(\regwritedata<0> ), .Y(n550) );
  AND2X2 U913 ( .A(n1036), .B(n832), .Y(n551) );
  INVX1 U914 ( .A(n551), .Y(n552) );
  AND2X2 U915 ( .A(n285), .B(\regwritedata<6> ), .Y(n553) );
  INVX1 U916 ( .A(n553), .Y(n554) );
  AND2X2 U917 ( .A(fow_EXID_rs_EX), .B(\regwritedata_m<12> ), .Y(n555) );
  INVX1 U918 ( .A(n555), .Y(n556) );
  AND2X2 U919 ( .A(fow_EXID_rs_EX), .B(\regwritedata_m<15> ), .Y(n557) );
  INVX1 U920 ( .A(n557), .Y(n558) );
  BUFX2 U921 ( .A(n1055), .Y(n559) );
  BUFX2 U922 ( .A(n1029), .Y(n560) );
  INVX1 U923 ( .A(n607), .Y(n561) );
  AND2X2 U924 ( .A(n285), .B(\regwritedata<2> ), .Y(n562) );
  INVX1 U925 ( .A(n562), .Y(n563) );
  INVX1 U926 ( .A(n880), .Y(n564) );
  AND2X2 U927 ( .A(n1036), .B(n660), .Y(n565) );
  INVX1 U928 ( .A(n565), .Y(n566) );
  AND2X1 U929 ( .A(\regwritedata_m<8> ), .B(fow_EXID_rt_EX), .Y(n567) );
  INVX1 U930 ( .A(n567), .Y(n568) );
  INVX1 U931 ( .A(n569), .Y(n570) );
  AND2X2 U932 ( .A(\regwritedata<4> ), .B(n1179), .Y(n571) );
  INVX1 U933 ( .A(n571), .Y(n572) );
  AND2X2 U934 ( .A(n1179), .B(\regwritedata<5> ), .Y(n573) );
  INVX1 U935 ( .A(n573), .Y(n574) );
  AND2X2 U936 ( .A(\regwritedata<6> ), .B(n1179), .Y(n575) );
  INVX1 U937 ( .A(n575), .Y(n576) );
  INVX1 U938 ( .A(n612), .Y(n577) );
  BUFX2 U939 ( .A(n1037), .Y(n578) );
  BUFX2 U940 ( .A(n1043), .Y(n579) );
  INVX1 U941 ( .A(n719), .Y(n580) );
  AND2X2 U942 ( .A(n191), .B(\forwarded_read2dataEX<12> ), .Y(n581) );
  INVX1 U943 ( .A(n581), .Y(n582) );
  AND2X2 U944 ( .A(\instIF_q<5> ), .B(n890), .Y(n583) );
  INVX1 U945 ( .A(n583), .Y(n584) );
  AND2X2 U946 ( .A(\instIF_q<14> ), .B(n890), .Y(n585) );
  INVX1 U947 ( .A(n585), .Y(n586) );
  AND2X2 U948 ( .A(\instIF_q<15> ), .B(n890), .Y(n587) );
  INVX1 U949 ( .A(n587), .Y(n588) );
  BUFX2 U950 ( .A(n1034), .Y(n589) );
  BUFX2 U951 ( .A(n1025), .Y(n590) );
  BUFX2 U952 ( .A(n1031), .Y(n591) );
  INVX1 U953 ( .A(n702), .Y(n592) );
  OR2X2 U954 ( .A(n1049), .B(n945), .Y(n702) );
  OR2X2 U955 ( .A(n1049), .B(n945), .Y(n593) );
  INVX1 U956 ( .A(n593), .Y(n594) );
  OR2X2 U957 ( .A(n308), .B(n965), .Y(n595) );
  INVX1 U958 ( .A(n595), .Y(n596) );
  AND2X2 U959 ( .A(\shamt<0> ), .B(n222), .Y(n597) );
  INVX1 U960 ( .A(n597), .Y(n598) );
  AND2X2 U961 ( .A(\immEX<0> ), .B(n925), .Y(n599) );
  INVX1 U962 ( .A(n599), .Y(n600) );
  AND2X2 U963 ( .A(n1045), .B(n861), .Y(n601) );
  INVX1 U964 ( .A(n601), .Y(n602) );
  INVX1 U965 ( .A(n603), .Y(n604) );
  INVX1 U966 ( .A(n605), .Y(n606) );
  AND2X2 U967 ( .A(\regwritedata<10> ), .B(n1179), .Y(n607) );
  AND2X2 U968 ( .A(n939), .B(n940), .Y(n608) );
  INVX1 U969 ( .A(n608), .Y(n609) );
  AND2X2 U970 ( .A(\regwritedata<9> ), .B(n285), .Y(n610) );
  INVX1 U971 ( .A(n610), .Y(n611) );
  AND2X2 U972 ( .A(\regwritedata<1> ), .B(n1179), .Y(n612) );
  INVX1 U973 ( .A(n612), .Y(n613) );
  BUFX2 U974 ( .A(n1021), .Y(n614) );
  INVX1 U975 ( .A(n615), .Y(n616) );
  BUFX2 U976 ( .A(n1177), .Y(n617) );
  INVX1 U977 ( .A(n621), .Y(n618) );
  AND2X2 U978 ( .A(n1020), .B(n837), .Y(n619) );
  INVX1 U979 ( .A(n619), .Y(n620) );
  AND2X2 U980 ( .A(\regwritedata<9> ), .B(n1179), .Y(n621) );
  OR2X2 U981 ( .A(n841), .B(n737), .Y(n622) );
  INVX1 U982 ( .A(n622), .Y(n623) );
  AND2X2 U983 ( .A(n222), .B(\shamt<3> ), .Y(n624) );
  INVX1 U984 ( .A(n624), .Y(n625) );
  INVX1 U985 ( .A(n547), .Y(n626) );
  OR2X2 U986 ( .A(n289), .B(n1014), .Y(n627) );
  INVX1 U987 ( .A(n627), .Y(n628) );
  AND2X2 U988 ( .A(n554), .B(n560), .Y(n629) );
  INVX1 U989 ( .A(n629), .Y(n630) );
  INVX1 U990 ( .A(n629), .Y(n631) );
  AND2X2 U991 ( .A(n802), .B(n305), .Y(n632) );
  AND2X2 U992 ( .A(n649), .B(n561), .Y(n634) );
  AND2X2 U993 ( .A(n546), .B(n576), .Y(n635) );
  INVX1 U994 ( .A(n635), .Y(n636) );
  INVX1 U995 ( .A(n635), .Y(n637) );
  AND2X2 U996 ( .A(n572), .B(n665), .Y(n638) );
  INVX1 U997 ( .A(n638), .Y(n640) );
  AND2X2 U998 ( .A(n552), .B(n1027), .Y(n641) );
  INVX1 U999 ( .A(n641), .Y(n642) );
  INVX1 U1000 ( .A(n641), .Y(n643) );
  AND2X2 U1001 ( .A(n725), .B(n568), .Y(n644) );
  INVX1 U1002 ( .A(n644), .Y(n645) );
  INVX1 U1003 ( .A(n644), .Y(n646) );
  AND2X2 U1004 ( .A(n727), .B(n570), .Y(n647) );
  INVX1 U1005 ( .A(n647), .Y(n648) );
  BUFX2 U1006 ( .A(n1182), .Y(n649) );
  BUFX2 U1007 ( .A(n1202), .Y(n650) );
  AND2X2 U1008 ( .A(fow_EXID_rt_EX), .B(\regwritedata_m<5> ), .Y(n651) );
  INVX1 U1009 ( .A(n651), .Y(n652) );
  BUFX2 U1010 ( .A(n1180), .Y(n653) );
  AND2X2 U1011 ( .A(\regwritedata<0> ), .B(n1179), .Y(n654) );
  INVX1 U1012 ( .A(n654), .Y(n655) );
  AND2X2 U1013 ( .A(fow_MEMID_rs_EX), .B(n1048), .Y(n656) );
  INVX1 U1014 ( .A(n656), .Y(n657) );
  INVX1 U1015 ( .A(n656), .Y(n658) );
  OR2X2 U1016 ( .A(n661), .B(n980), .Y(n659) );
  AND2X2 U1017 ( .A(n1011), .B(n189), .Y(n660) );
  AND2X2 U1018 ( .A(\regwritedata_m<14> ), .B(fow_EXID_rs_EX), .Y(n661) );
  INVX1 U1019 ( .A(n662), .Y(n663) );
  INVX1 U1020 ( .A(n803), .Y(n664) );
  INVX1 U1021 ( .A(n664), .Y(n665) );
  INVX1 U1022 ( .A(\regwritedata<5> ), .Y(n666) );
  INVX1 U1023 ( .A(n666), .Y(n667) );
  INVX1 U1024 ( .A(n301), .Y(n668) );
  INVX1 U1025 ( .A(n404), .Y(n669) );
  INVX1 U1026 ( .A(n646), .Y(n1191) );
  INVX1 U1027 ( .A(n285), .Y(n670) );
  INVX1 U1028 ( .A(jump_ID), .Y(n1183) );
  INVX1 U1029 ( .A(n671), .Y(n672) );
  INVX1 U1030 ( .A(n673), .Y(n674) );
  OR2X1 U1031 ( .A(n682), .B(n676), .Y(n675) );
  OR2X1 U1032 ( .A(n684), .B(n683), .Y(n676) );
  AND2X2 U1033 ( .A(n191), .B(fow_EXID_rt_EX), .Y(n677) );
  INVX1 U1034 ( .A(n677), .Y(n678) );
  INVX1 U1035 ( .A(\read2dataID<0> ), .Y(n1117) );
  INVX1 U1036 ( .A(\read2dataID<1> ), .Y(n1118) );
  INVX1 U1037 ( .A(\read2dataID<2> ), .Y(n1119) );
  INVX1 U1038 ( .A(\read2dataID<3> ), .Y(n1120) );
  INVX1 U1039 ( .A(\read2dataID<4> ), .Y(n1121) );
  INVX1 U1040 ( .A(\read2dataID<5> ), .Y(n1122) );
  INVX1 U1041 ( .A(\read2dataID<6> ), .Y(n1123) );
  INVX1 U1042 ( .A(\read2dataID<7> ), .Y(n1124) );
  INVX1 U1043 ( .A(\read2dataID<8> ), .Y(n1125) );
  INVX1 U1044 ( .A(\read2dataID<9> ), .Y(n1126) );
  INVX1 U1045 ( .A(\read2dataID<10> ), .Y(n1127) );
  INVX1 U1046 ( .A(\read2dataID<11> ), .Y(n1128) );
  INVX1 U1047 ( .A(\read2dataID<12> ), .Y(n1129) );
  INVX1 U1048 ( .A(\read2dataID<13> ), .Y(n1130) );
  INVX1 U1049 ( .A(\read2dataID<14> ), .Y(n1131) );
  INVX1 U1050 ( .A(\read2dataID<15> ), .Y(n1132) );
  INVX1 U1051 ( .A(\read1dataID<0> ), .Y(n1133) );
  INVX1 U1052 ( .A(\read1dataID<1> ), .Y(n1134) );
  INVX1 U1053 ( .A(\read1dataID<2> ), .Y(n1135) );
  INVX1 U1054 ( .A(\read1dataID<3> ), .Y(n1136) );
  INVX1 U1055 ( .A(\read1dataID<4> ), .Y(n1137) );
  INVX1 U1056 ( .A(\read1dataID<5> ), .Y(n1138) );
  INVX1 U1057 ( .A(\read1dataID<6> ), .Y(n1139) );
  INVX1 U1058 ( .A(\read1dataID<7> ), .Y(n1140) );
  INVX1 U1059 ( .A(\read1dataID<8> ), .Y(n1141) );
  INVX1 U1060 ( .A(\read1dataID<9> ), .Y(n1142) );
  INVX1 U1061 ( .A(\read1dataID<10> ), .Y(n1143) );
  INVX1 U1062 ( .A(\read1dataID<11> ), .Y(n1144) );
  INVX1 U1063 ( .A(\read1dataID<12> ), .Y(n1145) );
  INVX1 U1064 ( .A(\read1dataID<13> ), .Y(n1146) );
  INVX1 U1065 ( .A(\read1dataID<14> ), .Y(n1147) );
  INVX1 U1066 ( .A(\read1dataID<15> ), .Y(n1148) );
  AND2X1 U1067 ( .A(n1160), .B(n1005), .Y(n680) );
  INVX1 U1068 ( .A(n680), .Y(n681) );
  AND2X1 U1069 ( .A(\instIF_q<11> ), .B(n1178), .Y(n682) );
  AND2X1 U1070 ( .A(\instIF_normal<11> ), .B(n992), .Y(n683) );
  BUFX2 U1071 ( .A(n124), .Y(n992) );
  OR2X1 U1072 ( .A(jump_ID), .B(jump_EX), .Y(n684) );
  AND2X2 U1073 ( .A(\regwritedata_m<11> ), .B(fow_EXID_rt_EX), .Y(n685) );
  INVX1 U1074 ( .A(n685), .Y(n686) );
  INVX1 U1075 ( .A(n687), .Y(n688) );
  AND2X2 U1076 ( .A(n892), .B(fow_EXID_rt_EX), .Y(n689) );
  INVX1 U1077 ( .A(n689), .Y(n690) );
  INVX1 U1078 ( .A(n691), .Y(n692) );
  AND2X2 U1079 ( .A(n196), .B(fow_EXID_rt_EX), .Y(n693) );
  INVX1 U1080 ( .A(n693), .Y(n694) );
  BUFX2 U1081 ( .A(n1194), .Y(n695) );
  BUFX2 U1082 ( .A(n1195), .Y(n696) );
  BUFX2 U1083 ( .A(n1189), .Y(n697) );
  BUFX2 U1084 ( .A(n1190), .Y(n698) );
  BUFX2 U1085 ( .A(n1193), .Y(n699) );
  BUFX2 U1086 ( .A(n1198), .Y(n700) );
  BUFX2 U1087 ( .A(n1201), .Y(n701) );
  INVX1 U1088 ( .A(n702), .Y(n703) );
  AND2X1 U1089 ( .A(n974), .B(n1197), .Y(n704) );
  INVX1 U1090 ( .A(n704), .Y(n705) );
  INVX1 U1091 ( .A(n706), .Y(n707) );
  INVX1 U1092 ( .A(n1015), .Y(n708) );
  INVX1 U1093 ( .A(n708), .Y(n709) );
  INVX1 U1094 ( .A(n710), .Y(n711) );
  INVX1 U1095 ( .A(n712), .Y(n713) );
  INVX1 U1096 ( .A(n714), .Y(n715) );
  AND2X1 U1097 ( .A(n1045), .B(n835), .Y(n716) );
  INVX1 U1098 ( .A(n716), .Y(n717) );
  BUFX2 U1099 ( .A(n800), .Y(n718) );
  INVX1 U1100 ( .A(n891), .Y(n719) );
  AND2X1 U1101 ( .A(n953), .B(n954), .Y(n720) );
  INVX1 U1102 ( .A(n720), .Y(n721) );
  INVX1 U1103 ( .A(n722), .Y(n723) );
  AND2X1 U1104 ( .A(\read2dataEX<8> ), .B(n1042), .Y(n724) );
  INVX1 U1105 ( .A(n724), .Y(n725) );
  AND2X2 U1106 ( .A(\read2dataEX<13> ), .B(n1042), .Y(n726) );
  INVX1 U1107 ( .A(n726), .Y(n727) );
  AND2X1 U1108 ( .A(\read2dataEX<14> ), .B(n1042), .Y(n728) );
  INVX1 U1109 ( .A(n728), .Y(n729) );
  AND2X1 U1110 ( .A(instMemStall), .B(jump_IF), .Y(n730) );
  INVX1 U1111 ( .A(n730), .Y(n731) );
  AND2X1 U1112 ( .A(branch_if), .B(instMemStall), .Y(n732) );
  INVX1 U1113 ( .A(n732), .Y(n733) );
  AND2X1 U1114 ( .A(instMemDone_q), .B(\instIF_q<11> ), .Y(n734) );
  INVX1 U1115 ( .A(n734), .Y(n735) );
  AND2X1 U1116 ( .A(n1045), .B(n864), .Y(n736) );
  INVX1 U1117 ( .A(n736), .Y(n737) );
  INVX1 U1118 ( .A(n1041), .Y(n738) );
  AND2X1 U1119 ( .A(n877), .B(n858), .Y(n739) );
  INVX1 U1120 ( .A(n739), .Y(n740) );
  BUFX2 U1121 ( .A(n1033), .Y(n741) );
  INVX1 U1122 ( .A(n741), .Y(n968) );
  OR2X1 U1123 ( .A(DcacheErr), .B(IcacheErr), .Y(err) );
  INVX1 U1124 ( .A(n678), .Y(n1032) );
  AND2X1 U1125 ( .A(\read2dataEX<0> ), .B(n1042), .Y(n743) );
  AND2X1 U1126 ( .A(\read2dataEX<7> ), .B(n1042), .Y(n744) );
  AND2X1 U1127 ( .A(\read2dataEX<10> ), .B(n1042), .Y(n745) );
  BUFX2 U1128 ( .A(instMemDone_d), .Y(n746) );
  AND2X1 U1129 ( .A(n966), .B(n1197), .Y(n747) );
  INVX1 U1130 ( .A(n747), .Y(n748) );
  AND2X1 U1131 ( .A(\regwritedata_m<6> ), .B(fow_EXID_rt_EX), .Y(n749) );
  INVX1 U1132 ( .A(n749), .Y(n750) );
  AND2X1 U1133 ( .A(n983), .B(n1197), .Y(n751) );
  INVX1 U1134 ( .A(n751), .Y(n752) );
  INVX1 U1135 ( .A(n753), .Y(n754) );
  BUFX2 U1136 ( .A(n902), .Y(n755) );
  BUFX2 U1137 ( .A(\forwarded_read2dataEX<9> ), .Y(n756) );
  BUFX2 U1138 ( .A(n1206), .Y(n757) );
  BUFX2 U1139 ( .A(\forwarded_read2dataEX<5> ), .Y(n758) );
  BUFX2 U1140 ( .A(\forwarded_read2dataEX<4> ), .Y(n759) );
  INVX1 U1141 ( .A(n760), .Y(n761) );
  INVX1 U1142 ( .A(n762), .Y(n763) );
  INVX1 U1143 ( .A(n764), .Y(n765) );
  INVX1 U1144 ( .A(n766), .Y(n767) );
  INVX1 U1145 ( .A(n648), .Y(n1187) );
  INVX1 U1146 ( .A(n768), .Y(n769) );
  INVX1 U1147 ( .A(n770), .Y(n771) );
  INVX1 U1148 ( .A(n772), .Y(n773) );
  AND2X2 U1149 ( .A(n863), .B(n695), .Y(n774) );
  INVX1 U1150 ( .A(n774), .Y(n775) );
  AND2X2 U1151 ( .A(n861), .B(n696), .Y(n776) );
  INVX1 U1152 ( .A(n776), .Y(n777) );
  INVX1 U1153 ( .A(n778), .Y(n779) );
  INVX1 U1154 ( .A(n780), .Y(n781) );
  INVX1 U1155 ( .A(n782), .Y(n783) );
  INVX1 U1156 ( .A(n784), .Y(n785) );
  AND2X1 U1157 ( .A(\immEX<8> ), .B(n186), .Y(n786) );
  AND2X1 U1158 ( .A(\immEX<13> ), .B(n186), .Y(n787) );
  AND2X1 U1159 ( .A(\immEX<14> ), .B(n925), .Y(n788) );
  AND2X2 U1160 ( .A(n930), .B(fow_EXID_rt_EX), .Y(n789) );
  INVX1 U1161 ( .A(n789), .Y(n790) );
  AND2X1 U1162 ( .A(n931), .B(n1197), .Y(n791) );
  INVX1 U1163 ( .A(n791), .Y(n792) );
  AND2X1 U1164 ( .A(n973), .B(n1197), .Y(n793) );
  INVX1 U1165 ( .A(n793), .Y(n794) );
  INVX1 U1166 ( .A(\regwritedata_m<2> ), .Y(n1014) );
  BUFX2 U1167 ( .A(n1176), .Y(n795) );
  INVX1 U1168 ( .A(n795), .Y(n1178) );
  BUFX2 U1169 ( .A(memwrite), .Y(n796) );
  INVX1 U1170 ( .A(n297), .Y(n797) );
  OR2X1 U1171 ( .A(instMemDone_q), .B(n1203), .Y(n798) );
  INVX1 U1172 ( .A(n798), .Y(n799) );
  AOI22X1 U1173 ( .A(\immEX<7> ), .B(n186), .C(n285), .D(\regwritedata<7> ), 
        .Y(n800) );
  INVX1 U1174 ( .A(n1181), .Y(n801) );
  INVX1 U1175 ( .A(n801), .Y(n802) );
  AOI21X1 U1176 ( .A(\read1dataEX<4> ), .B(n1056), .C(n1050), .Y(n803) );
  INVX1 U1177 ( .A(n805), .Y(n804) );
  BUFX2 U1178 ( .A(n98), .Y(n805) );
  INVX1 U1179 ( .A(n807), .Y(n806) );
  BUFX2 U1180 ( .A(n83), .Y(n807) );
  INVX1 U1181 ( .A(n809), .Y(n808) );
  BUFX2 U1182 ( .A(n81), .Y(n809) );
  INVX1 U1183 ( .A(n811), .Y(n810) );
  BUFX2 U1184 ( .A(n79), .Y(n811) );
  INVX1 U1185 ( .A(n813), .Y(n812) );
  BUFX2 U1186 ( .A(n77), .Y(n813) );
  INVX1 U1187 ( .A(n815), .Y(n814) );
  BUFX2 U1188 ( .A(n75), .Y(n815) );
  INVX1 U1189 ( .A(n817), .Y(n816) );
  BUFX2 U1190 ( .A(n73), .Y(n817) );
  INVX1 U1191 ( .A(n819), .Y(n818) );
  BUFX2 U1192 ( .A(n71), .Y(n819) );
  INVX1 U1193 ( .A(n821), .Y(n820) );
  BUFX2 U1194 ( .A(n69), .Y(n821) );
  INVX1 U1195 ( .A(n823), .Y(n822) );
  BUFX2 U1196 ( .A(n65), .Y(n823) );
  INVX1 U1197 ( .A(n825), .Y(n824) );
  BUFX2 U1198 ( .A(n96), .Y(n825) );
  INVX1 U1199 ( .A(n827), .Y(n826) );
  BUFX2 U1200 ( .A(n91), .Y(n827) );
  INVX1 U1201 ( .A(n829), .Y(n828) );
  BUFX2 U1202 ( .A(n89), .Y(n829) );
  BUFX2 U1203 ( .A(n87), .Y(n830) );
  BUFX2 U1204 ( .A(n85), .Y(n831) );
  INVX1 U1205 ( .A(n833), .Y(n832) );
  AND2X2 U1206 ( .A(\immEX<5> ), .B(n186), .Y(n833) );
  AND2X1 U1207 ( .A(\read2dataEX<11> ), .B(n1042), .Y(n834) );
  INVX1 U1208 ( .A(n834), .Y(n835) );
  INVX1 U1209 ( .A(n1022), .Y(n836) );
  INVX1 U1210 ( .A(n836), .Y(n837) );
  INVX1 U1211 ( .A(n836), .Y(n838) );
  AND2X1 U1212 ( .A(\read1dataEX<13> ), .B(n1056), .Y(n839) );
  INVX1 U1213 ( .A(n839), .Y(n840) );
  INVX1 U1214 ( .A(n660), .Y(n841) );
  OR2X2 U1215 ( .A(n994), .B(n735), .Y(n842) );
  AND2X1 U1216 ( .A(\read2dataEX<4> ), .B(n1042), .Y(n843) );
  INVX1 U1217 ( .A(n843), .Y(n844) );
  AND2X1 U1218 ( .A(\read2dataEX<6> ), .B(n1042), .Y(n845) );
  INVX1 U1219 ( .A(n845), .Y(n846) );
  AND2X1 U1220 ( .A(\read2dataEX<9> ), .B(n1042), .Y(n847) );
  INVX1 U1221 ( .A(n847), .Y(n848) );
  INVX1 U1222 ( .A(n850), .Y(n849) );
  AND2X1 U1223 ( .A(\read2dataEX<5> ), .B(n1042), .Y(n850) );
  INVX1 U1224 ( .A(n851), .Y(n852) );
  BUFX2 U1225 ( .A(n223), .Y(n853) );
  BUFX2 U1226 ( .A(\opB<13> ), .Y(n854) );
  AND2X2 U1227 ( .A(n995), .B(n799), .Y(n855) );
  INVX1 U1228 ( .A(n855), .Y(n856) );
  INVX1 U1229 ( .A(n855), .Y(n857) );
  BUFX2 U1230 ( .A(n1199), .Y(n858) );
  BUFX2 U1231 ( .A(n655), .Y(n859) );
  AND2X1 U1232 ( .A(\read2dataEX<2> ), .B(n1042), .Y(n860) );
  INVX1 U1233 ( .A(n860), .Y(n861) );
  AND2X2 U1234 ( .A(\read2dataEX<3> ), .B(n1042), .Y(n862) );
  INVX1 U1235 ( .A(n862), .Y(n863) );
  INVX1 U1236 ( .A(n865), .Y(n864) );
  AND2X1 U1237 ( .A(\read2dataEX<1> ), .B(n1042), .Y(n865) );
  INVX1 U1238 ( .A(n867), .Y(n866) );
  AND2X1 U1239 ( .A(\read1dataEX<9> ), .B(n1056), .Y(n867) );
  INVX1 U1240 ( .A(n307), .Y(n869) );
  BUFX2 U1241 ( .A(n544), .Y(n871) );
  BUFX2 U1242 ( .A(n637), .Y(n874) );
  BUFX2 U1243 ( .A(n228), .Y(n875) );
  BUFX2 U1244 ( .A(n633), .Y(n876) );
  INVX1 U1245 ( .A(n878), .Y(n877) );
  AND2X2 U1246 ( .A(fow_MEMID_rt_EX), .B(n1045), .Y(n878) );
  INVX1 U1247 ( .A(n830), .Y(n8) );
  INVX1 U1248 ( .A(n831), .Y(n9) );
  INVX1 U1249 ( .A(\r_wr<0> ), .Y(n1165) );
  INVX1 U1250 ( .A(\r_wr<1> ), .Y(n1166) );
  INVX1 U1251 ( .A(\r_wr<2> ), .Y(n1167) );
  INVX1 U1252 ( .A(id_rd_v), .Y(n1096) );
  INVX1 U1253 ( .A(\immID<7> ), .Y(n1115) );
  INVX1 U1254 ( .A(\regwritedata_m<1> ), .Y(n1012) );
  BUFX2 U1255 ( .A(n908), .Y(n879) );
  AND2X2 U1256 ( .A(n913), .B(\shamt<1> ), .Y(n880) );
  INVX1 U1257 ( .A(n993), .Y(n883) );
  BUFX2 U1258 ( .A(\regwritedata_m<15> ), .Y(n881) );
  INVX1 U1259 ( .A(n979), .Y(n946) );
  INVX1 U1260 ( .A(n900), .Y(n1185) );
  AND2X2 U1261 ( .A(instMemDone_q), .B(n995), .Y(n918) );
  INVX1 U1262 ( .A(n995), .Y(n993) );
  INVX1 U1263 ( .A(n993), .Y(n884) );
  INVX8 U1264 ( .A(n1006), .Y(n885) );
  INVX8 U1265 ( .A(n1002), .Y(n886) );
  BUFX2 U1266 ( .A(\regwritedata<14> ), .Y(n887) );
  BUFX2 U1267 ( .A(\regwritedata<15> ), .Y(n888) );
  BUFX4 U1268 ( .A(n857), .Y(n889) );
  AOI21X1 U1269 ( .A(\read1dataEX<7> ), .B(n1056), .C(n1054), .Y(n891) );
  BUFX2 U1270 ( .A(\regwritedata_m<7> ), .Y(n892) );
  AND2X2 U1271 ( .A(\regwritedata_m<7> ), .B(fow_EXID_rs_EX), .Y(n1054) );
  AND2X2 U1272 ( .A(n558), .B(n899), .Y(n959) );
  INVX1 U1273 ( .A(\aluOut<1> ), .Y(n893) );
  INVX1 U1274 ( .A(n893), .Y(n894) );
  AND2X2 U1275 ( .A(\aluOut<3> ), .B(n886), .Y(\wr_aluOut<3> ) );
  INVX4 U1276 ( .A(n1006), .Y(n1001) );
  INVX4 U1277 ( .A(n1006), .Y(n1000) );
  INVX4 U1278 ( .A(n1006), .Y(n999) );
  BUFX2 U1279 ( .A(\instMEM_normal<12> ), .Y(n895) );
  INVX1 U1280 ( .A(\aluOut<4> ), .Y(n896) );
  INVX1 U1281 ( .A(n896), .Y(n897) );
  AND2X2 U1282 ( .A(\regwritedata<8> ), .B(n1179), .Y(n898) );
  OR2X1 U1283 ( .A(n1007), .B(n986), .Y(n900) );
  INVX1 U1284 ( .A(n1012), .Y(n901) );
  INVX1 U1285 ( .A(n975), .Y(n926) );
  BUFX2 U1286 ( .A(n962), .Y(n903) );
  NOR3X1 U1287 ( .A(n976), .B(n977), .C(n898), .Y(n904) );
  INVX1 U1288 ( .A(\regwritedata_m<3> ), .Y(n905) );
  INVX1 U1289 ( .A(n905), .Y(n906) );
  BUFX4 U1291 ( .A(n1205), .Y(n908) );
  INVX1 U1292 ( .A(n993), .Y(n1004) );
  BUFX2 U1293 ( .A(n213), .Y(n910) );
  INVX1 U1294 ( .A(n203), .Y(n911) );
  AND2X2 U1295 ( .A(n549), .B(n959), .Y(n970) );
  BUFX2 U1296 ( .A(\regwritedata<12> ), .Y(n912) );
  AND2X2 U1297 ( .A(shift), .B(n1036), .Y(n913) );
  INVX1 U1298 ( .A(n881), .Y(n1044) );
  AND2X2 U1299 ( .A(\aluOut<2> ), .B(n886), .Y(\wr_aluOut<2> ) );
  AND2X2 U1300 ( .A(\aluOut<10> ), .B(n886), .Y(\wr_aluOut<10> ) );
  AND2X2 U1301 ( .A(n958), .B(jump_ID), .Y(n1184) );
  AND2X2 U1302 ( .A(\aluOut<9> ), .B(n886), .Y(\wr_aluOut<9> ) );
  BUFX2 U1303 ( .A(rst), .Y(n914) );
  INVX1 U1304 ( .A(\aluOut<9> ), .Y(n915) );
  INVX1 U1305 ( .A(n915), .Y(n916) );
  INVX1 U1306 ( .A(instMemDone_q), .Y(n1204) );
  INVX1 U1307 ( .A(n1004), .Y(n1003) );
  BUFX2 U1308 ( .A(\instMEM_normal<14> ), .Y(n917) );
  INVX1 U1309 ( .A(\aluOut<12> ), .Y(n919) );
  INVX1 U1310 ( .A(n919), .Y(n920) );
  INVX1 U1311 ( .A(n1014), .Y(n921) );
  AND2X1 U1312 ( .A(n922), .B(\immEX<3> ), .Y(n924) );
  INVX1 U1313 ( .A(n191), .Y(n922) );
  INVX1 U1314 ( .A(shift), .Y(n923) );
  AND2X2 U1315 ( .A(n922), .B(n923), .Y(n925) );
  BUFX2 U1316 ( .A(\instWB_normal<15> ), .Y(n927) );
  BUFX2 U1317 ( .A(\instMEM_normal<13> ), .Y(n928) );
  INVX1 U1318 ( .A(n224), .Y(n929) );
  INVX1 U1319 ( .A(n797), .Y(n1186) );
  BUFX2 U1320 ( .A(\regwritedata_m<9> ), .Y(n930) );
  BUFX2 U1321 ( .A(\regwritedata<6> ), .Y(n931) );
  BUFX2 U1322 ( .A(n928), .Y(n932) );
  BUFX2 U1323 ( .A(\aluOut<10> ), .Y(n933) );
  INVX1 U1324 ( .A(\aluOut<5> ), .Y(n934) );
  INVX1 U1325 ( .A(n934), .Y(n935) );
  AND2X2 U1326 ( .A(n563), .B(n1018), .Y(n936) );
  BUFX2 U1327 ( .A(n912), .Y(n937) );
  BUFX2 U1328 ( .A(\aluOut<13> ), .Y(n938) );
  INVX1 U1329 ( .A(n670), .Y(n939) );
  INVX1 U1330 ( .A(n1026), .Y(n940) );
  INVX1 U1331 ( .A(\regwritedata<4> ), .Y(n1026) );
  BUFX2 U1332 ( .A(\instMEM_normal<11> ), .Y(n941) );
  INVX1 U1333 ( .A(\instWB_normal<12> ), .Y(n942) );
  INVX1 U1334 ( .A(n942), .Y(n943) );
  BUFX2 U1335 ( .A(n906), .Y(n944) );
  AND2X1 U1336 ( .A(\read1dataEX<0> ), .B(n1056), .Y(n945) );
  INVX4 U1337 ( .A(n995), .Y(n994) );
  INVX1 U1338 ( .A(n979), .Y(n947) );
  AND2X1 U1339 ( .A(\read1dataEX<14> ), .B(n1056), .Y(n980) );
  INVX4 U1340 ( .A(n963), .Y(\forwarded_read1dataEX<12> ) );
  INVX1 U1341 ( .A(n182), .Y(n948) );
  BUFX2 U1342 ( .A(\instWB_normal<13> ), .Y(n949) );
  BUFX2 U1343 ( .A(n870), .Y(n950) );
  AND2X2 U1344 ( .A(\aluOut<15> ), .B(n886), .Y(\wr_aluOut<15> ) );
  BUFX2 U1345 ( .A(\instWB_normal<14> ), .Y(n951) );
  BUFX2 U1346 ( .A(\instMEM_normal<15> ), .Y(n952) );
  INVX1 U1347 ( .A(n1036), .Y(n953) );
  INVX1 U1348 ( .A(n1035), .Y(n954) );
  INVX1 U1349 ( .A(\aluOut<11> ), .Y(n955) );
  INVX1 U1350 ( .A(n955), .Y(n956) );
  BUFX2 U1351 ( .A(n895), .Y(n957) );
  INVX1 U1352 ( .A(br_ctl), .Y(n958) );
  BUFX2 U1353 ( .A(n888), .Y(n960) );
  AND2X2 U1354 ( .A(n650), .B(n577), .Y(n961) );
  AND2X2 U1355 ( .A(n559), .B(n556), .Y(n963) );
  BUFX2 U1356 ( .A(\regwritedata<10> ), .Y(n964) );
  AND2X2 U1357 ( .A(\read1dataEX<11> ), .B(n1056), .Y(n965) );
  BUFX2 U1358 ( .A(\regwritedata<9> ), .Y(n966) );
  NOR3X1 U1359 ( .A(n679), .B(n968), .C(n969), .Y(n967) );
  AND2X2 U1360 ( .A(\read1dataEX<15> ), .B(n1056), .Y(n971) );
  BUFX2 U1361 ( .A(\regwritedata<3> ), .Y(n972) );
  INVX4 U1362 ( .A(n1174), .Y(n995) );
  INVX1 U1363 ( .A(n212), .Y(n1192) );
  BUFX2 U1364 ( .A(n667), .Y(n973) );
  BUFX2 U1365 ( .A(n887), .Y(n974) );
  NOR3X1 U1366 ( .A(n977), .B(n976), .C(n978), .Y(n975) );
  AND2X2 U1367 ( .A(fow_EXID_rs_EX), .B(\regwritedata_m<8> ), .Y(n976) );
  AND2X2 U1368 ( .A(\read1dataEX<8> ), .B(n1056), .Y(n977) );
  AND2X2 U1369 ( .A(\regwritedata<8> ), .B(n1179), .Y(n978) );
  NOR3X1 U1370 ( .A(n661), .B(n980), .C(n981), .Y(n979) );
  AND2X2 U1371 ( .A(\regwritedata<14> ), .B(n1179), .Y(n981) );
  BUFX2 U1372 ( .A(\regwritedata<0> ), .Y(n982) );
  INVX1 U1373 ( .A(n1026), .Y(n983) );
  AND2X2 U1374 ( .A(n545), .B(n574), .Y(n984) );
  BUFX4 U1375 ( .A(n914), .Y(n985) );
  BUFX4 U1376 ( .A(rst), .Y(n986) );
  INVX8 U1377 ( .A(n987), .Y(n988) );
  INVX8 U1378 ( .A(n987), .Y(n989) );
  INVX4 U1379 ( .A(n877), .Y(n1197) );
  INVX4 U1380 ( .A(n1008), .Y(n1042) );
  INVX4 U1381 ( .A(n657), .Y(n1179) );
  BUFX4 U1382 ( .A(n856), .Y(n990) );
  INVX8 U1383 ( .A(n1005), .Y(n996) );
  INVX8 U1384 ( .A(n1005), .Y(n997) );
  INVX8 U1385 ( .A(n994), .Y(n1005) );
  INVX2 U1386 ( .A(fow_EXID_rt_EX), .Y(n1045) );
  OR2X2 U1387 ( .A(fow_EXID_rt_EX), .B(fow_MEMID_rt_EX), .Y(n1008) );
  OR2X2 U1388 ( .A(n193), .B(n1009), .Y(n1010) );
  OR2X2 U1389 ( .A(shift), .B(n1010), .Y(n1011) );
  OAI21X1 U1390 ( .A(n1045), .B(n1012), .C(n219), .Y(n1013) );
  AOI21X1 U1391 ( .A(n623), .B(n225), .C(n616), .Y(n1207) );
  AND2X2 U1392 ( .A(\shamt<2> ), .B(n222), .Y(n1017) );
  NAND3X1 U1393 ( .A(\immEX<2> ), .B(n923), .C(n1036), .Y(n1015) );
  OAI21X1 U1394 ( .A(n289), .B(n861), .C(n709), .Y(n1016) );
  NOR3X1 U1395 ( .A(n1016), .B(n628), .C(n1017), .Y(n1018) );
  AOI21X1 U1396 ( .A(n1045), .B(n863), .C(n1019), .Y(n1022) );
  NAND3X1 U1397 ( .A(n620), .B(n785), .C(n625), .Y(n1021) );
  AOI21X1 U1398 ( .A(n838), .B(n906), .C(n614), .Y(n1023) );
  OAI21X1 U1399 ( .A(n844), .B(n208), .C(n711), .Y(n1024) );
  AOI21X1 U1400 ( .A(n191), .B(n851), .C(n1024), .Y(n1025) );
  OAI21X1 U1401 ( .A(n846), .B(n1036), .C(n713), .Y(n1028) );
  AOI21X1 U1402 ( .A(\regwritedata_m<6> ), .B(n1032), .C(n1028), .Y(n1029) );
  OAI21X1 U1403 ( .A(n848), .B(n1036), .C(n715), .Y(n1030) );
  AOI21X1 U1404 ( .A(\regwritedata_m<9> ), .B(n1032), .C(n1030), .Y(n1031) );
  AOI22X1 U1405 ( .A(\immEX<10> ), .B(n186), .C(n191), .D(n745), .Y(n1033) );
  OAI21X1 U1406 ( .A(n1188), .B(\regwritedata_m<11> ), .C(n717), .Y(n1035) );
  AOI22X1 U1407 ( .A(\immEX<11> ), .B(n186), .C(n285), .D(\regwritedata<11> ), 
        .Y(n1034) );
  AOI22X1 U1408 ( .A(\read2dataEX<12> ), .B(n1042), .C(n912), .D(n1197), .Y(
        n1037) );
  OAI21X1 U1409 ( .A(n1045), .B(n1038), .C(n578), .Y(
        \forwarded_read2dataEX<12> ) );
  OAI21X1 U1410 ( .A(n1047), .B(n1039), .C(n582), .Y(\opB<12> ) );
  NAND3X1 U1411 ( .A(n191), .B(n1197), .C(\regwritedata<13> ), .Y(n1040) );
  NAND3X1 U1412 ( .A(n191), .B(n1197), .C(n887), .Y(n1041) );
  AOI22X1 U1413 ( .A(\read2dataEX<15> ), .B(n1042), .C(n888), .D(n1197), .Y(
        n1043) );
  OAI21X1 U1414 ( .A(n1045), .B(n1044), .C(n579), .Y(
        \forwarded_read2dataEX<15> ) );
  OAI21X1 U1415 ( .A(n1047), .B(n1046), .C(n300), .Y(\opB<15> ) );
  OR2X2 U1416 ( .A(fow_EXID_rs_EX), .B(fow_MEMID_rs_EX), .Y(n1053) );
  AND2X2 U1417 ( .A(n196), .B(fow_EXID_rs_EX), .Y(n1049) );
  AOI22X1 U1418 ( .A(fow_EXID_rs_EX), .B(n901), .C(\read1dataEX<1> ), .D(n1056), .Y(n1202) );
  AOI22X1 U1419 ( .A(fow_EXID_rs_EX), .B(n921), .C(\read1dataEX<2> ), .D(n1056), .Y(n1180) );
  AOI22X1 U1420 ( .A(fow_EXID_rs_EX), .B(\regwritedata_m<3> ), .C(
        \read1dataEX<3> ), .D(n1056), .Y(n1181) );
  AOI22X1 U1421 ( .A(\read1dataEX<5> ), .B(n1056), .C(n184), .D(fow_EXID_rs_EX), .Y(n1051) );
  AOI22X1 U1422 ( .A(\read1dataEX<6> ), .B(n1056), .C(fow_EXID_rs_EX), .D(
        \regwritedata_m<6> ), .Y(n1052) );
  NAND3X1 U1423 ( .A(n618), .B(n866), .C(n869), .Y(\forwarded_read1dataEX<9> )
         );
  AOI22X1 U1424 ( .A(fow_EXID_rs_EX), .B(\regwritedata_m<10> ), .C(
        \read1dataEX<10> ), .D(n1056), .Y(n1182) );
  AOI22X1 U1425 ( .A(\read1dataEX<12> ), .B(n1056), .C(n1179), .D(
        \regwritedata<12> ), .Y(n1055) );
  NAND3X1 U1426 ( .A(n310), .B(n626), .C(n840), .Y(\forwarded_read1dataEX<13> ) );
  OR2X2 U1427 ( .A(br_ctl), .B(haltMEM), .Y(n1174) );
  AND2X2 U1428 ( .A(\aluOut<0> ), .B(n886), .Y(\wr_aluOut<0> ) );
  AND2X2 U1429 ( .A(\aluOut<1> ), .B(n886), .Y(\wr_aluOut<1> ) );
  AND2X2 U1430 ( .A(\aluOut<4> ), .B(n1005), .Y(\wr_aluOut<4> ) );
  AND2X2 U1431 ( .A(\aluOut<5> ), .B(n1005), .Y(\wr_aluOut<5> ) );
  AND2X2 U1432 ( .A(\aluOut<6> ), .B(n1005), .Y(\wr_aluOut<6> ) );
  AND2X2 U1433 ( .A(\aluOut<7> ), .B(n1005), .Y(\wr_aluOut<7> ) );
  AND2X2 U1434 ( .A(\aluOut<8> ), .B(n1005), .Y(\wr_aluOut<8> ) );
  AND2X2 U1435 ( .A(\aluOut<11> ), .B(n886), .Y(\wr_aluOut<11> ) );
  AND2X2 U1436 ( .A(\aluOut<12> ), .B(n886), .Y(\wr_aluOut<12> ) );
  AND2X2 U1437 ( .A(\aluOut<13> ), .B(n886), .Y(\wr_aluOut<13> ) );
  AND2X2 U1438 ( .A(\aluOut<14> ), .B(n886), .Y(\wr_aluOut<14> ) );
  NAND3X1 U1439 ( .A(n1175), .B(instMemDone_q), .C(n1183), .Y(n1176) );
  AOI22X1 U1440 ( .A(\instIF_normal<0> ), .B(n991), .C(\instIF_q<0> ), .D(
        n1178), .Y(n98) );
  OAI21X1 U1441 ( .A(n805), .B(n889), .C(n520), .Y(\wr_instIF<0> ) );
  AOI22X1 U1442 ( .A(\instIF_normal<1> ), .B(n991), .C(\instIF_q<1> ), .D(
        n1178), .Y(n83) );
  OAI21X1 U1443 ( .A(n807), .B(n889), .C(n522), .Y(\wr_instIF<1> ) );
  AOI22X1 U1444 ( .A(\instIF_normal<2> ), .B(n991), .C(\instIF_q<2> ), .D(
        n1178), .Y(n81) );
  OAI21X1 U1445 ( .A(n809), .B(n990), .C(n524), .Y(\wr_instIF<2> ) );
  AOI22X1 U1446 ( .A(\instIF_normal<3> ), .B(n991), .C(\instIF_q<3> ), .D(
        n1178), .Y(n79) );
  OAI21X1 U1447 ( .A(n811), .B(n889), .C(n526), .Y(\wr_instIF<3> ) );
  AOI22X1 U1448 ( .A(\instIF_normal<4> ), .B(n991), .C(\instIF_q<4> ), .D(
        n1178), .Y(n77) );
  OAI21X1 U1449 ( .A(n813), .B(n990), .C(n528), .Y(\wr_instIF<4> ) );
  AOI22X1 U1450 ( .A(\instIF_normal<5> ), .B(n991), .C(\instIF_q<5> ), .D(
        n1178), .Y(n75) );
  OAI21X1 U1451 ( .A(n815), .B(n990), .C(n584), .Y(\wr_instIF<5> ) );
  AOI22X1 U1452 ( .A(\instIF_normal<6> ), .B(n991), .C(\instIF_q<6> ), .D(
        n1178), .Y(n73) );
  OAI21X1 U1453 ( .A(n817), .B(n889), .C(n530), .Y(\wr_instIF<6> ) );
  AOI22X1 U1454 ( .A(\instIF_normal<7> ), .B(n991), .C(\instIF_q<7> ), .D(
        n1178), .Y(n71) );
  OAI21X1 U1455 ( .A(n819), .B(n990), .C(n532), .Y(\wr_instIF<7> ) );
  AOI22X1 U1456 ( .A(\instIF_normal<8> ), .B(n992), .C(\instIF_q<8> ), .D(
        n1178), .Y(n69) );
  OAI21X1 U1457 ( .A(n821), .B(n889), .C(n534), .Y(\wr_instIF<8> ) );
  AOI22X1 U1458 ( .A(\instIF_normal<9> ), .B(n992), .C(\instIF_q<9> ), .D(
        n1178), .Y(n65) );
  OAI21X1 U1459 ( .A(n823), .B(n990), .C(n536), .Y(\wr_instIF<9> ) );
  AOI22X1 U1460 ( .A(\instIF_normal<10> ), .B(n992), .C(\instIF_q<10> ), .D(
        n1178), .Y(n96) );
  OAI21X1 U1461 ( .A(n825), .B(n990), .C(n538), .Y(\wr_instIF<10> ) );
  AOI22X1 U1462 ( .A(n1203), .B(n1204), .C(n675), .D(n855), .Y(n1177) );
  NAND3X1 U1463 ( .A(n617), .B(n842), .C(n1004), .Y(\wr_instIF<11> ) );
  AOI22X1 U1464 ( .A(\instIF_normal<12> ), .B(n992), .C(\instIF_q<12> ), .D(
        n1178), .Y(n91) );
  OAI21X1 U1465 ( .A(n827), .B(n889), .C(n540), .Y(\wr_instIF<12> ) );
  AOI22X1 U1466 ( .A(\instIF_normal<13> ), .B(n992), .C(\instIF_q<13> ), .D(
        n1178), .Y(n89) );
  OAI21X1 U1467 ( .A(n829), .B(n889), .C(n542), .Y(\wr_instIF<13> ) );
  AOI22X1 U1468 ( .A(\instIF_normal<14> ), .B(n992), .C(\instIF_q<14> ), .D(
        n1178), .Y(n87) );
  OAI21X1 U1469 ( .A(n830), .B(n990), .C(n586), .Y(\wr_instIF<14> ) );
  AOI22X1 U1470 ( .A(\instIF_normal<15> ), .B(n992), .C(\instIF_q<15> ), .D(
        n1178), .Y(n85) );
  OAI21X1 U1471 ( .A(n831), .B(n990), .C(n588), .Y(\wr_instIF<15> ) );
  OAI21X1 U1472 ( .A(n203), .B(n658), .C(n580), .Y(n1205) );
  NOR3X1 U1473 ( .A(jump_IF), .B(n1185), .C(n1184), .Y(pc_en) );
  AOI21X1 U1474 ( .A(n909), .B(n1197), .C(n1188), .Y(n1189) );
  AOI21X1 U1475 ( .A(n964), .B(n1197), .C(n745), .Y(n1190) );
  NAND3X1 U1476 ( .A(n848), .B(n748), .C(n790), .Y(\forwarded_read2dataEX<9> )
         );
  OAI21X1 U1477 ( .A(n877), .B(n1192), .C(n1191), .Y(
        \forwarded_read2dataEX<8> ) );
  AOI21X1 U1478 ( .A(n197), .B(n1197), .C(n744), .Y(n1193) );
  NAND3X1 U1479 ( .A(n846), .B(n750), .C(n792), .Y(n1206) );
  NAND3X1 U1480 ( .A(n849), .B(n652), .C(n794), .Y(\forwarded_read2dataEX<5> )
         );
  NAND3X1 U1481 ( .A(n844), .B(n752), .C(n852), .Y(\forwarded_read2dataEX<4> )
         );
  AOI22X1 U1482 ( .A(n972), .B(n1197), .C(n944), .D(fow_EXID_rt_EX), .Y(n1194)
         );
  AOI22X1 U1483 ( .A(n948), .B(fow_EXID_rt_EX), .C(n231), .D(n1197), .Y(n1195)
         );
  AOI21X1 U1484 ( .A(n929), .B(fow_EXID_rt_EX), .C(n1196), .Y(n1199) );
  AOI21X1 U1485 ( .A(n982), .B(n1197), .C(n743), .Y(n1198) );
  NAND3X1 U1486 ( .A(n740), .B(n754), .C(n191), .Y(n1201) );
endmodule

